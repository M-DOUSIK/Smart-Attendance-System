PK   x#X�i%X,  X�    cirkitFile.json���Ʊ�_e����FF^x�o�maؖ`�|���R�����n�dA�/�ϴ��U�ؕ���h�;[�ӕ�����Ŷ�g�j7�~��~{���\��py�C����/k./ޭoVw������o�gw?��f��]��Ǭב	ݐٺ�3ߕ!����
�*WOe�Vfe.�~����Hl��H� �`VV� �`VN� �`V^� �`VA� �`V��Aj��
1�ԂY�b����R1G���D� �Jy�$y����t)6)�	Sl"R�S��D��'M��H!O�b�B�8�&"�<u�Mı�<w�MD
y������<wZy�����)6)�Sl"R�s��D���N��H!ϝb�B�;�&�&��N��H!ϝb�B�;�&"@��s���N��H!ϝb�B�;�&"�<w�MD
y�M<h7?����7w��0u��*+��e>EV��gC^y(��*r�@�wG��m���l[���V�6��v}�sv�/�"/��b�B���&"�<��MD
y����Vy��.6)�9\l"R�s�h���YJs�<��MD
y�0� ϻb�B�w�&"�<�&Ώ�B�A���&"�<g�MD
�#2y��-6)�9[l"R���D���]�	���yWl"R���D���݉��z�<˙w�ۙ4^t��˲�LQי�|�Jg�O}�����P��������]M/fNNg�A ݞ9��t��3+�����JGX:�rX߹C����e�^M/L�'�u�ǆ,���tq��]��JGX�8���.��JGX:�*��+�����άJ��J��t��3�
�
�;(a��]L�,J�|��H��C�2Kk�,����]����x����9��4�|�㷥���,���=o�����G`>~C�?������߭��<�|��U`������|��<7�X>��J�����G`>^C�����XX���`���#0����?�|��G`������|�V
�?������Wy���X>���4�����G`>^Y�X`���k��w�����|���?�������a���X>��
R�����G`>^�
�X`��ǫv���,��x�1�`���#0����?�|��5�`������|���!�����x]�.�|�^��],_<X�`�������,����`���#0O �,_�|��`����W�����/X>�q������G`>.�X�`���%J���,����
���'X>�qY��X`���m���,����`���#0��?�|��F`������|\|	������s}_���B�YcL�{7d5ue64����v������FG.M�*�t	`��#0���,]�|��*_`������|\����T'-D��gzi8{�"!`Փ�U���|\N�?�������t��R�^��� 9%\S���M��狋쮪}���2_�[u��LU�����ݸ��ٞ��J�OM�S[��ZV��HN�D�$�>�I��� "/$�����S�J}��3'|Xu��e�$]|��ݖ�s����l_��t-@	@��-*��`^x�a�䅇V=^x�a��=Aړ�]i�������ğv�a�����rp�mKr�}rW�SW�S��<vnT�8���znT�8���znT�8D��z�vy�~N���doĥ�ύ�
˾�B�� �Rxz/+ٹ�4='r�d�¥��ߔ�ec�ù@�L�I�ćIB/��j�2��}$&��1w#H,�.��.��\i�жY��|�����r�u��vh�W�g���NW��&�<^I�B��ˆ�u���~��I�ϟ���z�퐙�,3o���Y��]o�5�_9{�ᯜ}h}nJ���ƑD��e㳦)�����T��=�������:����UC��c��MF��d���(8�Ϟt�x�_��Ww�U���l/��r�-�0�������Rr�2|�"�!�yC2dxC2dxbC2dx~C2dx�C2dx�	C2dx2C2dx~C2d�)7P��em\چ�m�%n�%3N7��`��`�eɌӢ &X�&XGY2��-�	��	��Q��8�b��q��(Kf�"1��߸8,�[XGY2�L3�	��-,��,�qF�����Q��8b��q��(Kf�m�qXw�<���e�`L���T
,�;XGY�e0&Xw�<��ĥ�`L�<�`y��R�5A���;KTV����0aye�k��`y���8����1���q��<�aye����`y�����%
^��`ye�k_��`�� ��(K\������w�*�L��`ye���ØpO7q�7ay<��8�/��1�����Q���;,��<��īNaL�<�����%�����C���3�t�l�jV����V�~�`%V�:\F�
��+���3��aA�c�?g��V����Op��x�`%�8R��a'�4XI�5�QT�zX�	�VRa5��zOp�@�j��
�Yց�[�U��TX����*Я������ťBK:��n��o�T�����]�#�HGy�В-�k��[EC:��C�����VG��В-����[�BK:���AǷ:JL��thy-��ouԘ
-�����(2Zҡ�1:��Qe*��C�k|t,��2Zҡ�J:���e*��C�k�t|��DL鑘�.�:����2Zҡ�5p:���e*��C�k�t|���ThI���$��VG��В-����.S�%Z^#��[]�BK:���UǷ:�L��thyͮ΋I:�L��thy�out�
-���j���2Zҡ��:���e*��C�k�u|���ThI������VG��В-���.S�%Z����[]�BK:�\�AǷ:�L��th�v��o�J��AG��E8���2���ThI��k���VG��В-�D��.S�%Z���[]�BK:�\�FǷJ+ɔ����2��˼�.S�%Z���[]�BK:�\�HǷ:�L��th����out�
-��r-*��</S�%Z����۠��ThI��k���VG��В-�8��.S�%Z�զ�[]�BK:�\sNǷ:�L��th���D�v�t�*�t��]tt�
-��r-C���2Zҡ嚌:���e*��C;���-�`��eGh�f�u�ttY���ThI��k}��VG��В-�,U�	�T� �`Gh!�M�e/�/rWվ͊�w��ݐU��3SU>/ꢰC�ۇ�
ƸZ`e�M;�+z���j�ap���۱��X�������je���I`e�n]�Ɣ���Q�1yq��P��qy�U�2�"+}�!/�<]O3�o�B+3��Z��>�Њ���OI���h���j����/_he���B+35F(x1�;�I�R3c�d�K33�;�R3�~أ����f�<u�L3S��3�e=s�6�f��=;͌=usJ3�Ň;�-5��⹽C��y�⺗�x���n)K�<��Í����8�K����.&��6�l��m7�Pe66�|�F5ue64����v��w�����IV�g���Sc���}^�mf���<�CV:���7}�:���$+t*������ʕ�m����̷����,�]�!o��==�L�r:^\i�j����B�f�]6�������i�$+'Y������i�2󦡬nj��}����ZC�4K���,C�sS�,�6j�<D+e㳦)�xA�k��+'Y��u�ol���!�n�z��MF��d���(�O�$Yy���hfu�Y���w���_��.߆��n���m}��o�., Cf�VȐ3�dȌjB2dF�	!2�����QC�@�̨�!D CfT�"�!3�~Ȑ�� `R$.k��6,o,q�,��D	�	��	��Q��n
���K�(Kf7��a��p�%q�%����0���q�%����0��߸8,�[XGY2�yG,�[XGY2�Q,�[XGY2��Z,�[XGY2�Yd���q��(K\�Ƅ�I�M����q�%��c��q��(K\������Q��n�	��=,��,q�,�{XGY�0&ܜ8nR��=,��,q�,�{XGY���0&X��<����a�~`y<��8���1��x��q�%^
c�=��=ބ�� ��(K�N�����Q�x]�	��sXGY�uP0&X�ay|���5M�5sh���G ���J*�f5Y/��
��+����d��*Я���jV��%h�@�j��
k�]*~��.�x@��TX�8Hů��%h��
k���uR��VRa5�I��U�_5XI�լ&�J�V�~�`%V���)A[�U��TX��`a���ThI���m���R�]:��t��(/Zҡ�w�u|���ThI��ߙ��S�%Z~�_Ƿ:*L��thy��ou��
-���Z��1Zҡ�5%:��Qd*��C�kct|���ThI�����<X��e*��C�k�t|���ThI���\��V鉘�#1]fut���e*��C�k�t|���ThI������VG��В-�I��.S�%Z^[��[]�BK:��FTǷ:�L��thy���out�
-���]��tt�
-����c���2Zҡ�5�:���e*��C�k�u|������:����2���ThI������VG��В-���.S�%Z����[]�BK:�\�AǷ:�L��th�v��out�
-��r�z]�BK:�\KDǷ:�L��th�&��out�
-��rm���2Zҡ�5:�UZI���LG�y]�ut�
-��r� ���2Zҡ��G:���e*��C�5�t|���ThI��kQ��VG��В-��R�m��e*��C˵�t|���ThI��k���VG��В-�j��.S�%Z�9��[]�BK:�\;OǷJU>��|�負�˂�.S�%Z�e��[]�BK:�\�QǷ:�L��th����out�
-��r�L��:�L��th�֧�out�
-��r�R���2ZJ�}��x����mV���|톬�|����yQ���}�Z��M���L5مVf�x/�2Sy{���Z���T�^he�����0u��*+��e>EV��gC^y(�*��t�$Y9/IVN�K����d�d�$Y9/IVN�K�L��T_he�F�Ҩ/&z�6	^j�s[�.5���o�����ܶ�K�`�xn�֥f@9�s��.5��⹽C���D���K�`�xn̥w]L��6�l��m7�Pe���>��j��lhr[��\ݟ�$Y����PE���,��u�yʇ�t6�ԗ�o��u8}EIVN^Q����zW�>�mB�3��>+C(��w]h���6A��X9���P�6Y?�Q��*d�лl(<9_]��xI�r����z�퐙�,3o���Y��]o�5�O�$Y9�2�>7��Bk���C�R6>k������T	,)VN���:���%WC���rk��o�4��Q*�dI�������Ow�vs�ٮ��Oo�^^�_o��ջ����f��v����7�<����۠o�|w���I6`�n�P��@�6l��W(E�ѴxJD2m 9s.rKN���Jrj'SO�S[�⒜�Ȥ���$�{�>k+S�\�>���BzzW���9)N)��l�K�W�k�!�����D�&B18+�Ԥ�A����S%A��ٛU��M:}�ݣ(��?n�UI}�(�D������KU�T�ǿ�T<B���������~�忉?������QD��x��C����r霁�@:u '�� �	�	r�|`�V�P�g �I�t���H�M��o��Ή��o2�*�o1%"όȿ3���H:O"����%<a����f��������O������n��_wo��}~*�zɻ<��M�񩶐Bl�)�&�����Bl�)�&�����Bl�/)�&�����Bl�O)�&�����Bl���ߖ�-D�D�O@�$@��0�WХ�J�$*�av/�K9 y� �Tn��^×r r)��܆�-�r ��S��[� �@�GR@>��|*�av�)��|j�Tn���sH9 ���܆٭(�r ��S��[�"���|� �Tn�w	p >B���S�ީ�ȧ�O�6x  �:@>m��?d�X��:�8�"�d[��� �ȶ�m�6�N>�1���Rd[ȶr\��ȶ�mG���TB,@����� �`6 ҫ��%p �k �����]�� �Vn�+�8O��� �6 ���W�p ƶ�^�6��  ���*��o8 �5�ש�+D�t-|=yRyR�KS\�= �YM�L��A���#0�YM
I��A���#0��x�M����z
��Wx����8{�p���/�>����^/���|q� �ߤ��z�|�3�I�}�=���|�3�I}�=���|�3�I�|�=���|��7 ��i� ����D�.J�-K�K-L���&�f�>Ď�	MHhB~��C�"���VF��J���&�7��>D+0!�	�-q���LHhB~��C�B����G��R���&��yk�N��WE�}��)`BB���P�OP�:Ţu�E�0!�	y%ڇh�&$4!�B��S���&�Lh�u
��Є��
�C�N��W��}��)`BB�7��:LHhB^��~?�S���&�Նh�u
��Є�R�C�N��Wy�}��)`BB�
U��:LHhB^]��!Z��		M�+��>D�0!�	yU3ڇh�&$4!��F��S���&�/1���D�����e�X���--[���&�e�h�e��Є\r �C�l���%�}��-`BBr���S�+Sвţe�G�0!�	��ڇh�&$4!�A�-[���&���C�l��밠}�~�&$4!א�0�u
��Є\��C�N��k��}��)`BBr�!��:LHhB.���!Z��		M���Ƈp0��= _T��--[Z��		M�u��>D�0!�	�Fڇh�&$4�tS�I6s8���U��K���2G�0!�	�XBb|�V1`���֓
����ͼ'�E�s�~��_�8�wW�\��FÉ[%O��슛�����̶���iO����dnR�u���/0�O������Ĝd��I�Υ[y��T�\��=��D"[h�H(I�M���]x��t���'%o?)U�4���*���K8��W�[��IA��aHGr�L�M�7�fd�n�fo�?��)-�����/���������ܢ��M�2I��t۶��!o�7qy|�Hrc�Gz@%�wd�I��n$���+�;ic�i��O�g>�?I�l�0� ���?r�3�5qK���O2w�b����}h�,��g��}V�Pf���y;��k#ؤ�_�,W��&�<J�P��z��'���}�������]_�Cm�̴e�y�PV7���>�zSWm�^_;��h}nJ���FA��x|���i�:���5ի�O9������:����UC���wk��o�4��Qu�r���w�������u��۬��ۋ��\�Ȳ���\pg���:�-��8��'�]^�d�ӆ./��qvo����uLhcG�ӘAƬ4�V�#,aG�|��#,a��GX>����p|D̾?%���ǃR2�䠔~�|�%t��Rz��	��w@J�ퟡ���)B6�E<���CSeM&oj��[���!㐉�[�UDydiB�lev-���n�mִ���&��l롯��o�]��Z��綪زn��616]շщC�kY�j�2�}�r��d�5}�|�:��k��M�Zj���r�P��"��ǀa�UݵƆ�j���2+��g6ƁsM�G܇+�u�K
Y쁑3~'�{��Ѹ��s!ܮ�-�.PQgUUƖ��Ř���*bǋ�ִv�=�~��o�;�����)��` ::�#	�p�é�)���K���Ma�F$��/���R*��	�D2ƻӔ&�Ј�9BSHh$�.޾�4��F2�i�M�Gs��"�;!"#$
��9ҷ��D����ÅSB+%M���4��%?��)�\�N��":s
n.�'JtY�����̞8Y}�nJ7��g�D�nS��L�8u#��|18���[]G�^�� ���k�����z���ه���#��~�>�ӏ��Ga�Q��Q>��x���~T>|TN?�>�&ѣ7h�zr�����:�BS�УGh�zt	M}B�>��S��)4�
=z%�㣾�]��^��6�����mR���ʮ�k{{6����;�6�z���;��e��W�ͻ~{��y�'^R̨���&6�(ث2Tyn.�����W��x��h���OjƱUU�*�]�I�**��貲�;[��um�������iw�$M.]^l��H]�.���_��m{�?\G�4�*\�>}�U�?_�/�7��,]���ǐ7�A>^��A���/�1v4N�vEy�Gag�*��^W�o)��_��i��x��X�}}w߭7ﷷ;o�]��G�ˋ���_�Ŗ�w�����w7���o������=���|������:��E������/o��^����>~x�o���]7�������_o����Ř��c}s?�����߾���mw��� H���V�S/�zY��W�ʗ�l]�o\VĈ�
oڬ6�������x{�Is�	�lg"�W�>�7�,�>rf�(G�1�ϴs6��/�=�f��6�]�oo���73��Mk������`���t�M�XK%�4[M?qn�?{L>{L1{L5w�3s�8�#�h3W&5�0~�6����Vաߏ�:cG�MC�h�I�m5	�����u��$����o'TVí��������7�=/}[�Sa.�CP�n����'���>7}f�=$�M�gU�E���R�S��J�y�2/M��?cL�1���"�c�v�r�էȁEN��ݖ��$�H@IO SF�!/�"h~4���F�o<����*sEn?��l���x9
YEyU<%��қpUX����˸)mW8�(k���\�)/�lL_R��v����,�!t�H�ܿgU����T�#W���H�<a|{�����!2O�1�le��hO�M�;�]ֆPg��7�������}gh(���*�=���a�&P���^�����o׻Kx�u�{���w����7o�O_����_���{�\w�o�����2����!*DSU�Ӎ���4�ۼ�y�yn�0�?ص�ث��Q������5�l�?������#q5	������7_o>�o��W�۾�܃���&�t���(�C��-lLv!�YS�.3�/b&�g��������0~�^�9��qrm��Dn���l9h/��>���cX��7� J�)/l���u4zw��\�a�B�����w���	�p����"��O�^�;\岦jCV6��Z盌\A�s�޹n/V���K�mS��m��<�܄��@����\�|}�-���������Ư�����?��o�m�7u�E����ۻ�{��?}7��͋��z�_ď�7���޾��ݼy���|������I�=>�}���'��y`�w�^���<\�������W����w?|�t��H���?��n�o�?l�7/;�3�a�g�n��~�χ��n����I[=��^5�Oh�ٟ?}A��ש�������G�>}��hNZ������H�7�߿���+�W���<T����%����Ua��W��Q1����kWUY�;�
�,���=�h3L�+)��������n��������ގꘟ:�혹/���2X��K��U�S�;�&�O�3����c�N�����1?u�ߠcFEW�JlY����=�^�7�����⎙��#ꘟ���_����?���)�WE�}�r�L�s�@t�Y�Ʌ���ä%^Q?���s�}ꇟ��쇶
W�%g(��<W�K�+~�\�˝��b����#��o���S_��?p_t���Pc��0e��+VW�,B��)���]1i��G����|��>�P?���)��x��Z"
9]���F���w�8f���֘R	�#������|ꑟz䇽?���BY9�#z^���������Tm�#ꍟ=���?u�{s��NH�B銒������+�x�B�(�ZO��J�Ȼc��� ؽ���}�x����*����ۋ,��݊�{���~`��WQ!�~�����M����:+��tx��{�Wۺ���W����翯����?��˷1aĀ���������g�ۋ�oc������|э�]�g4��tGL������������ޟq�m�1��w?�����o/x=��W���cb��߾���ˋ�_�[�h��+R���h3�Y���f�c�|U,o������[}����ߏ��??ƫW�ט����5��wi�:������a�3��xT��XZ�<?lu<����V��H\Z�+=����Yt��`��j��ӷ9iƫ�n�hf�"(��9��7����k�ӛMz��zc��9.j��m���q�_�a6n�����JmV�3��3Z���_�u��V.�oz�ք�׆������İ�<��a�I^|Sce�#a{�,�cQL㑊I�MhV���ݻE'��	ȱ���V�a;}0��8l6l��K����l{�l&��Oʶ͊�� ��/n5�UR�Vg��1ap2l-p�`�ak�a���8l�jK��㣾I����l?�Қ�=�G���n�&i�`�$p� W#�� �m	[�Ͷ�yak���l��7+��f����Vs��H	��Vɷ��PE��H�@#l~�������Yn&_�a��u�c��ar<ݪ�Gǘ� �&���z6�~�*��N��>�N�i`؞̏�|��}��ߧs���=+[������p|���L��V�7R�Lۀ�% ǀ'���,:X���no�5,�f&p����V������Ч2����'��D�`��)��U�#9c��	� (������^���YG(�d��V�?�S���&���h%$�i�Yc�EςӶ=�f��]҇�X�y���0�������9h5`~?��J}x�(t������93r�#��R}���s�l�~��s��Ϣw�����v�|ej*rx#ݼ����*����f3�/e�r��[N��RGK��'mO�M+�=X�7�#�KoZ�u��k�s�j&*�<%v[%���vޜ5�����-2X���_.`���z~��%4����}H���,�oL�'ρ���|��F~�mn�����%���)����A~Ik5j�������/�]�]�׷o9�n����w�o����6?~q��x���ů�PK   0�"X�l��z� S� /   images/02fd9929-a358-4090-8e7d-8cad28564328.png  @߿�PNG

   IHDR  �  +   ��u   sRGB ���   gAMA  ���a   	pHYs  �  ����e  ��IDATx^��׏eK���Y���Z߸ZeVʪʪlvO��� �!�	�o�Ð �db�C`�/6��Kk��:��U��.�="�}�ev�q�q3���n���mbٲe�~&��]��՗7��o�o�i�WW[۽��l�m=޶��b�oq�|��|���Y�;��ݻ����˶�i�m��/̷��Ŷ�������]�	�����&�677�Ƴg�~��⛅t��Li���e��}�;y쒞]�py����w��f��sо����y���w[�����iɍ\˚v,w��R4�yŚ�])k��U�W�}i�͙^ϟt��{Y���:���\�R$�/�!���s�}Z��i��Ԙ�N�|H�U�^e*q:)ڪ��a��z��x��r��<���"_�3�3��[��b���^&��"��H��.�q�K~ÚO�n��ӥ6�k.�)/�#��/��e�Q<�����f�I�0�u�/����re��Z�<(3?7ߖ�o9M��g�������y��T(���Է!�݈�̐�v+_���2Vd��>���&v7��G���Yi�c��'r��� �n��g섩)S�� /��"�K�$���&�$�n���Gx�KX~��g��s��R^u�.x"_�m�Z}��^܌��<O��\�）��a��@_0�/�.��7���{�y��<��N��Ћ�K����Nr�<S�]�:uJ����ȕ�/�q�����ͤ4�.�C��i��i+[Io��ϑ�q?�(~�Fn��a,�)�xW�]]���q�������?��O��j*��\��!G���Ӽ<3*�v_�z´�"\��)m��N�ț���(ʱ>��3�
���ݴa�Fy�t�T���_P�?-9�(��66�G�EF"��5~��ʤ��^ط,,��mc6�&��]Z^��h�yc����l)�	������h}X��2��~����]��:����m"C8�E��e&Ϸ���LBo�2�Y��̲?�8X%bHU���x������n�#w������ID��{��i�1���S���4(eGI�7�K�E]N�cY�{�|Sg�VZB���"�xo�~IS7	�
ǧӔ uU&�	�D.�]���웖����AK�]��7?}y���v��v����l�4_�(�(R ��E�����o��o	>��
�����h�6Z�	� \�-��@A�#�}�������S���b>\xʏLR!�r�\�-&��K�(�h��d��$.�r���t�ָՑT���6��o��W���	�H'��y�/7���/�N)j�Z3���'�1K���Oe���������=ɒgsXٜ��b���>[_G^6"7d����V@;�{���[���z��*ݪʧU^b�k��U�:��-�d1vf��n�S~�e;�Yc��t4��2n��(se�h�bd\��T����E�� �������K�m��dY���a
�Nsl�5�+�c�Y��K�5g��O���G����>N�*�8�Y�6�n
���������<�6^�j�*��?��?�|��� �ʜ�AO�cv��F�bK��5�^ 3�ޒ0iN�+|q��u6����C��
����ͮ/u���m����v;eT�U��O�F~�u����z&��Q��P�\��v����	c�9@` H�U��We?1����`G �(I�U��Է^\k+dpU��hz�8�p'�q��	�W��k���NJ�-�q;���S��m�f�$�T�����D4SG\��M)�7wQ��'�U�L�_"�e��b���:Z[_e���LnF>��|��������^p�+�2c�i ە�LZi�kk����	�d�ҶK�zev�UFn)�s�˲Go�?[g8����]zz�%�Tf�9t7�'��J����#��C,'&U�x�?Me�u�o91��w�uc���c�˅ޚ���wA
����$D�OݏpՆ�y�b3X���w�Sȳr��7��6�MZ%�ZS(���6p��������u�">��,r��6z��ݿw��ۻ���,�]�տ����^��>��J�}�Q{��-����a`m\c��e&�g��'s	��9�0�L�p6�g� �W�&T�x�Q�`�1,�(���M!��ِ�2�:�^Jl|�ʨ����줭���H��Ҙ?=}�:���xIW��$��F^��3�3si��6`����@��'�lZ	;�{<ߞ��5&ϺW�{�_n"�0�`3�{l:+�*�g(�5�avn��n�]y�����H�L�ׅ��S2 _��]yP��K^b{���z��O�LPf�<G����|9ö����mq��L8����D>'���|4�y��&iK��:������o]����g��L��[�u�򒸙�6>�>�;hF��2���z��G�h�_��&�z���O-&�Wi��{�I��YO��]�I䈎�zBW��pi��1�?z��-�,�=�M��T��i�3w�h���а�/՗䧄��z2�]pkַ��η�n$���M�+�����zKy��!bC�Kr]`e�ЕD�	�'?���阰i�d_&u+$7������C��5qRc����NR��ލQ�7�l�|��^nS6kb�Z��~�p>3@�!�g=/<�I���T�-������'��q��$��^�Ys������LS��O۳-����"��/\�'�N��L��U0��(g�{֘���Rl��>��]#�g�ن�B<ui�h����.�)�T��g�/z�{�%�2m|�x	3�wj&���	2��IH�#z�M|�h&q�:��^\y#���Hc�ES�r��D�����/&f�6k�E�&���X�5���G��g�EMd���p�]Ň�UOʐH%Y�>����g����g��[��Ѧy���ff<荬�Z�,/�lW��}+�Ё�m��_���O/ n/^mw<i�w/��P������m`ED���e$z/�Uí�K1��oa�qo�Q��hH`���~5�4\3|�|�3�ɳd�u��k�bdi�D�L+ojȑ��$\�p���t�����c^�T��)�̣�cf���ܺ�ͬ"B+ȵl�����cO�u���l«�הw�m�c�d���q�(�u�y�*�.���i�\�癝��姱g�m:
3��<(�jg$��U��`[�4��KWJ�IZ�U&�K��]L�]�$XN~ːK������0_0&�����0>�/*&A�"�Y9�k��Z �� R�e��rH��	?��y>6
M�v*&��W/�	�C<�ڟn�.�~��!�� �I�j�k��V��.6a���uֺ��O��BwY�_�k�0�����}8:�X�l���O[�R�1�1ސ��G��$�2��H�G��k~�Opl��qj�K���F�ȱzG�q]���5a�n~��xN��^C�u ����\�����[4��0�W�mOZ$���
3��83|ts�Tc=5wď��,�"NM�C�n'���w�ʙmN���q6�-PF�P�������������X��º��TU_%���;۩u=�2%ݔ���-m"��4u��j߂��z��5[�J�9Y���0�,���΢���j6['S���\���-�d[������F[}���������%;֔r�۳5�ȡ�tzc��� �f�;K���yE��w��Č��ц˫\n'�}6�a0o�j�2��.��-c���0�\]�>3���/�j�Hc$z�-�zP���ׄ�X��c_0zu�8�e��#�2%o����g�uk�XÔ^F������wp�� ��#ڮ����}�	���K�ڽ�����E�� #jEIR�0>���;��I1$?�RnL��V-Q~6�4����◙m��R���Fuk�QX6+�O��}NO�ܦ9}\B�I	��+����y\�W�6��h�����n��͎�/3��(���=	f�6���1�3�^a�;�nb�."_i��<�h�Q
Z_�I��#x�Bh��D��miq>{Jaa��J�;�"���<y��-#ʪ쳼�+Y�!��Ј+��v�ц��p4<�	�����2�w\t����T��h̫�'�0�c��rfV�,��ŵôӶӳ[�1=���K��$+�-��n�e󑃱D����,c�0�ʽ}������%�\�G�����uB����˴�	�X��`�����4MO�I
�����ğ�by�'M;Z��5c?��yN'�Y����	;�O�͟t��!���Z�q� N0��	��(Fs��/֤Be%����� `c�ԫ�(����T:m�c���9I:��?�W�"#Å��F�n˘W����?ƫg	��p{��ǭq�#����d��Đ:�a��'����1a���5��3��E�����D���l'I}�G�Jg҄�?��6I��`�l@.�k<۲ ����W�F�3�L@�66u�bT�I��{/��z3�a�a�(���n�A��,,��c��U��<��l�XEm��9�W�*�x�ܔ�%�ɳ�O�"�ҙv7�w��67�����^a(\�랕t�v1���bj�mx��z�q&b��nH���
�����6c]�N��������<�t�_����`�F�u�:���m����f�j��L�1����#��b�>7]����pt����Cٽ+�ȡ�m׿�/���O/^o.�h�����������(!T��X��c-�x�g33I��^IR��K ;ڍ ����2;s�a����ϧ�z�)Z���ҏk���>h�뺛��^������`F�AZ�H��w�o��@	�	��f�������d��L����u�0�ɶk�Ex��Nc�~Yf�]�Ly^��K�����77 �]GP_������J;|�@;tp;x`o[��y)7*Osr������t�V�
���-ť�iʁ3��?R�3�Me�ggU�w u�0U�<SYy���}>逺B�ҁG�f�Ho��M�I���ub�Eܺ��ӽM+mq�-��'�W�y���2���.Rl�r�_�$)��������<9q�]s����kf�tD��vo��О���gt	^�L��_ҍ���4�Y��i�S�o�M���	���Y�N�C����k�� ��^�k����&E�����j+��է�'�y[� f�X[[�|8���
IL.�Z>����liHyf����pS�`��;6	T�;�ȡ��@�Ք!����V:��s-رpI����1��I�n��%-_��'���I�nKK�'@�^?��˹�.O�$��7�EV�6���{�V�0n�u�wņ%�A�&�r5U%�ڱ3�ʹ�,H׌q�K�Y���=�(3(�6�$��7F��߆p�*T�q�;L���z'e��������]`�v�{nz�$6{97�mgV�0�q+;�������n�����Z��I��`F��J��gʫ�nL3��'�1��m�w�{���m��P�|X&� >V�	�	�3�S:i��l�dx$Ef��t��M?�xݎ摟i��ԥ})��]�{���/3�w��eq�<�h&��,��ER������oϢ��w^~z	p{�f��p�m���9�rF�h
_/H2�仓�Ƀ�I����ڬ�B�5�����xӱT弊)���TA��u�-
cD��E�A���No�8k5�3��ad⏴��]��v�����2vT�+M�r��Ӥ43����eQfg ����K�N�*�_��+�	Q�ۭ�5 ���z[\����N�<�^;w�X;rx_[^ZD�S�(�9�m:Ed�:��&�+\;�-:!;��?lh��s]��[c�e�=��r��BDƌbr�)eS�ɮ�������_.����1�-S��S��2�n�W��}�J�#�ī���ZoHC�\�� ��jF��	�x���%?�'V:� D�uC/)��`( � �+���^%��2Rֺ"����i.ۖ����2i�e6>�>���ғ}������֭�� |��yt6��Ty�E{�M��.�`kb���3wI[Z\FV�=z�2��Y	@1��cɧ@�u\<s���ڶ\~Ό����r��.�@n�cH�Q�j�� ��1�n�o}�Q��rQ�x���)G�Q�֝2�!�5�^���j ��/v�3����$#�k\y��$|�����am�)�rn	�W�>ǵ>u�(��G¹�]�<��겾���ܓId���/K��Q��6	�̩\�UF+������R�<����k�Ƞ�5�K/Jwd[可4�wd�x�n~~1��A����/�f_�'��mu�Y[_w�8��^��d:��hN��������
���f�e��Ĕ�4���Ռ;m��J~��?:��)C�q�t*�01z%l\��<���(����n:��0����$�4<��󿻉o�矿�0��5�����z�鹔+���t�p����Ӝ��R73��~�|A���c��FWe7�ܮ�m���_�����g��ڽ�� w�����6�kM���S���l�RjϷ�[�l)HBY����Q��A;M* ���Y;�H���������~��S�+{�)y�M���Z�L�*z���U��>/3�i����S��:�yU���$���_M��א
\��>�*p�[��Ξlo��Z���w�'��Y[fG���HbL���M(
o�%���?�����{b�b����t��Tf�P7<��2{=L��#�'����p��3�Їd:�Ճ�r{��]MC�N������+|uA#r��e�m���'!����ҥ�=��<9�F���^[���
C���>1�ǰ�W�&���vp[a&/��pK�Kr*�<�2�������-�qEO�Boѭ��o6��n���[q*ˡ��)��e*��R���<*��LC��H���O���Ôe�͕�D(of[+�u8��4C;�8����ৣQ��3\����*�t�I�f�Gݧ|��y�~iU�Z���`���Z�u,z�n����N�a�Ǌ�!�N��EG�'ua,�	SRp���*\�-�c�8��d�w��� ��k����O^��;�����ŵ��i^l\Zj���%|��<�(�oqz�&ݝ�ƅ?�Y=�g�5<W���p���M=�u�*cuҒm������ݹ��ݹ�ݹ��=}� �o߳��L�v�7+3uQΗ��݄��M:)?�&Iݔ���1#?\i���iy�#i�&���㾻��3q���	;Kf\~l7��dK��ϓ����e�`S�z���]��.1F����TJ��F�C��LL"��o�Ϲ�y��g�k�CGl7�� оg�ڼ������g[��+�[ߴTA����8��A\[yu��}�`\F�$�2�,��z!�A{a��3��a���F�t�{�6lY�H����y����~9��%�04fȋ���U�1Mc��i�r��l�ٰ\��"u��Iȟ~�3��2ӟc���j�3�)9�س����}�ie��������z�}��wڷ�����k���}����{
��js��QZ�>|� luv7���X�X�_$7!�����s;͡�� ��;5;�i�nF^�x7�?hf��u*�{�ܙLc��=��;{��$���5�?��$?&��[��`��d��HS�<$��Q 0M�䯀��.6�̗���5^��)�ĕ�O	g��&x�n3l�?����Ԝ�B��1[��_���գ��y�����i�2ޏ����u�5��0�3"u��_�Ą�{~�̰�Y���{cc�=x��jy���ۛ��tjT�ky%�t%Ic:�$��
�<_p��-��$�"Cs�����ɥ̶gZ"�����	�M�����S��E��Gf"�ݠGZ������v�Ɍ(e���z"�uAĄ���yh��Fi5'�:˟��O0�2�$~�p���J�<�N�|'���CO7�@�||���-,��y����_�]�T'e��³
]��5L��Ӥ�:I�ґOXe.G�e �r����j�r�n�|�f����v��c�˹�SfLO���q��&4�B�7�L|F�<�rX���Awm+��τ��I6����xmwG��n�;.�TR�����%�����([��*�����X�]�k�0�u��Li{�=|ڬ+7�)?G�tf�4���"̸yPf"�ez�1E�}M���]�	���?���gno n� t�[d��i!ͪVIV;3�n�tO%P�+;��2z&���a��Ym7N
��{��Q�u�_���+��&��*��0=/���Ҹ���Oe�V��_�3�õ�����0�p߽�<#m~vFÄ�_�S~�����x��L�|U��J#=
�Kq�5ac�I;rpo�����׿�A��o5���������'����Q��?s6)���>I|��A6/y�;��Q���
Te��=�]���N#g��G�s�l�۰esg�\{�S��a�6��y�.*ɘ��$��S�v\�]���]��1��G�TѶ]��,����W�I��ҸX�=O�ΙXg�rn1�&�����iL��p�cq�g1��Wϊ^�[^�巇��p���K7Ǩu:qS�0mfD��u'�y�nu5��{�.W���Kܪ�n,L\�UW\�.t��?�!�2^m���zD���4�؛�2K.�C$�Uޚ�Xw�>
����٨$�ַ���?OTm�0�`L�+k��ú���|�?��<UY�����vG�u^�Sוc���2��+'X�Yg��V� ��!,����@��ɖ�o�E�xRi:tc�0�qCg
�}�I�aD��ڼ�n��ٓ��#�m�vgZ*�������Z�a,�R����"`ҋ+ߋWc0��<�=��O�gn�_��r�ɏ?m7n�e�e,_�D_�Wz�fGFbF�������v�S>ÿh���af��ew���LCO��=IS���u�ۃ�w��;���b�~b��15ʟr�h���2l���	E�fȫ�=��ǒ�����;�c�a\�#����"��������d;�5��ɔ��>dfb�{_���ۊK��ڮ��!���.^�p��[����8�_73��j�3}<���IL���naX��w&6q���oӜ�Î��[*$lA1��2V���(C��Bt~�e�QqU��t��~?1�K_7�b[��23�õ��;�V��� �W�C��<�U���A�����^�[F~������ȡ}�׾�^���?h����N�8�<��2�����v��mb	n���'���4�Bn�e�]Q��,D>ֻ�S�1\�pT�e��mL�����W 9��y#�]���z����]&�K�r�<��*��`m��˄�<*���x���y�P�C��:}�^8��3�����^H�B�r�n�L'����{�c� 2��v��Bn��z̸���i�_ns�?�s`r%��U=�NQ/En�O����pC���z=xZ���6I/!���=hI�[����V�<�x]���J���wWZt��o]�[7a����,��^p�__�,pˣ����e��#6��2�F<��b	N;�)XNNφ>�\�:�kSLzz�뜀�I�+� E�O�k�O�T�/qm��M�i�i��JIwjB�6�2�O`V��5�y@.pိ!�2�l��i��;]&�zۇ��$�Y��U������@dvei>�r�8��l�=Y{�V�m����n"�ݚ������]O}���N�r�ϖ)n�M���f~e��3�'��9�X��{�h�}�ٍ���\h���ewm�9��kK���k|m�.3�n"cuQ�ČȘ�/�w���3Io��8�y�S��|u�\x1��!�܎�8%��~��G��j��q^e���<�1R���&�I^�Y~��;�d�V)��>����~]���lg�'q+�i���7M���Vc�qsW��O�~b�u�-=7�s�������������
�ڒb�S%����j4P��4v;�/d�1NOg��$���7-�0���4	��w����Ŕ�M��gi������2E���f�,W���'Yy8M�ٞ�0�	���HJ���l3�H^Z�#���L����_b�����m"�i��0���n�8���������o}�>x�ݿ�%�Q�����O/��&������/2<�����Gkaz�7�(�T��n~w	j����	�L�f�JCD����'(���׆11���
�'�Ug7����3�;#_誣\f�-n���h�}q�@NeY�D�{�&ݢ������S�x�y%=c�I3��y�"?��[�-�q���@��g��+J����b�ޛj�d���%4�
I�h�g�t2�<�ۊW&�C\��7!���8�e�V����s@�&U?�����AG�9S���+q���X����$��g���iO�~mz��4wYN�愍<̼@�A�Y�-�Y{��a�?t�P��L�h�,�J��D^0��Zn��޼�r�n�%���M�@��M��iB��/�y�s)a��4���}�ز�E6ґ���*b����緗~vy�q�\c���������nd�� ���~�C��N�&��F� ���=��]T�ms���/�Sz�gj���v���n��-WF]��w���>Ў=@���U*�ӷ��mw>j�V}	�y�_��(���`����g��/taӾb{�1������
3�	�2*/꿤IQ)��2`|Ϟ����v����_ep�م[��?�����.\��V�nR�Wo�r\Oclq��*/MdK�:��\��Li���f�5̶tƣ�lR��wWã�у���~#�u1�[��wboG�֠	�#�+Ml;�+���,	�l��ť��Z|-Z�u�b�G��~�
���T��x�|r3���r]m�[~�ɥ�3�q�]�C���+��e����^>�p������vL��[?z(0����`$(�>���K�4p��%�\�c�ag�G�_��LN���;��{g����7�W�a�Ň��<0ĩx��?+>%��_af�wS��bG�$�����=L�o�4ّ�T9t�{2I|�׶��Ds�3r�/3�x�@J�JAod�vo��7��A�ַ~�ط7KZ��������;�>��s��me߁��R���H���ֲ�����@�ܼkg.8���PϾ�Ig�Z9��N	𻋎HP�K�ħΠ�t(Oo�m}��z���.0������Rօ���l�Q%L��K�[��}nQ7�̯��g�n�p<�M�%�6��k�	��T���`{SR?<�~i;�,Y;�^��tko�%!]�,�	����~����|��o�-;:Z�a"�7��k�a�9p�|���/4>�K�^�����^��[�K&�d-,��o�r�$b;�7N�7ס�k&�2�O��x��U��̤�-��|+ϕ�ʪ �3����O���?�����l����# �3JMY0�!���F��[Jx�ג������Ť-"�r�c��Z�e����lErP��d[O�O�Hډ�|8!vb3�t���� �)��D(_R4i���\>�Я?܎	����e�����/
�b����h��/�)��� 2A��A���S|ym���o��-���>t`O;s�h{�����[����J�{�i�v�N���v��v��h�bp�>j���Sx�̜(�ra��3�t9�&�eA��2T���C����>�/������Џ�]��� �#ǎ��gN���<���>�x��p��������ړ'�uw[;�kK6�R�p���N�W�n�n��;�0�C���g�L��:�5���"��45K.�G7O��7���u�GL�ʝЀ�|���6����Ы|��h�x���e�d	w)uo����(�>��@n�'�_F�<Ueq��*�n��ʉ�����f^T��Ck���Y^Ξ��@jY�	�'q8f/6v�>��`�k���U|�0�������Q?�my�,p�������ǟ_hx���:v�ȏ��7x)�}6k"X6f��a�������U%t4�a5~jf�G���M�ZW��ݬ�f62~�q�ͯ��u�1k���d^�Vaz���R���lbBH]v3���j�_�6n����m�g�2��1%w����O�)S�N���ف�`�����W�n_���׿�ݿ������������_\���h�)8��]�q��V��X��M�M b��/���,/eyv�8KX'�N���h� [mum�=y�wcï�I7���]��{����ZX�<G�Q��N����	ۑɃx���<hƹ�s���`�N����͊���#X�c	� �E�ޡI������ۓյ���@�@�7uy�� 6�Q�̂3�x*�&Q�=B�`-/.�M��
����`����*�ulRN딼Q��,�yJ�3R�v1��R�x����{�Ie�BPಥt�Y��U!���������iK���� ����Í�FJ_'o��s�9�S�[~q�<����A�nǐ��*�䅴�3��ݻ����m$������>O�O�_���K�����G��y�M�U�b4�B���f8'^f�,9*�8�������<��<�"�@���٭,���"��qNu�uQ �<(g� ��2M|M���?�:����,B?��󭍒�&�M��yFy���t�C�����6���_eR�� "2����]�A�'M)�ϥW�8������1K@N��nɳi�9�RVݲI��������2Q^iW�2{.�)V�A��m`���'t[���emj�{yw���v������l������{�K�O>�P�y��ҥv��m�ʳ� <?�G"�F�3�y[.�f��L dg�C��UY��4��Mk`��[g�.��+)�&�Z/�[6/����Ok��v���~��e@�9t�����_��On=\�@|qe�+p[ ��qꎟI߇[~�
a|&��6���`��^$t��6�c��%�Ȁu��!�=d\�Y�V� ��O���ޮ�����I' �Ȉ������3{m���ږҞ�X������'O�h'ObOO�'�}�.��>y�=�� {�=�w�m�����ߙ�gڑ#��2ịK�'rد�����O��0غ���א�����S�5V��++S��8���ӧb��w�m^S�X��5�����m���P{���N����p{��}�I�x)n�Z9��J��^m*G��*A	_��J�_�M�WH��F��?��Rش�Y�ý��xf>�2����L�H���͸����r��$������f6�\���I�hf��z���U��(հ_a����&�=�m�H��|��\[���>��и#3��6I�B�����h�����f��O����﷏?��b�+p{�H��MIA��� k�.���:}��� ����{i�ؽ{��={2�]���֞��3��f�<Ym�<̊���k 0?}j�EW�yt���AcVn�yt�f�5����pfn��kX�۽���;�k�����v9{%������]*��Yr�fP�tu�=B�<�}���:�o�CwΖt��E'+vTae��6k����+�^D�hW�������
���]x��s��x�� h�����)�
�EP�������#x�B��:|g`!���(`��-��q����P�L�a� �U��>�O�e' ݙ���6z[_D��sf��e�T\f^��+v�\��Fx�g�y�(�|m�m<\0�z����R�ч�33�;� bɁt
:�$��>tb-μo/Y+���j�:{�����׋����JڃKٖ�9�/&��:���s�*�d�%��DV�?� �*B?u���hXP,bs>���^J���mr��*l�d�5��a��-K��,���%'��|��gB孠`�Mڭ#�}Fy�m�z��$�~P�-`m?'�pBϯ[�"�*8-ms�.���	
�y=_�TT�m��ZpC.��Y�s������a+r ߵ�fd+`�2�CW���O�o~���O��w����ڧ�j?���������g��wn�7ۡ����}���_t�c�H��X������WxȀ:�ԁ�EGZ;���m�ve/t��l�c6�S��3A?|ܻO;y�D��7?l��_��v�رvAp��K�o����9v�� �w^pK�pk�-3�~5�M>�&R��<��C�1��>�C'E^1���s����^��]�k&��Hy��`�U�j�gz��	����8U�}��-�ȇp�;��ef���IwQB�n���V���v������~��?��;{
�� �I߶��}��q�u�V�q�z�z�J{��q����c���o�N����{��ZQp�k��oܼ�.^��ce�1�����w�����mX�g�'O��}�}�n� +3�"*iO�2[������I���En���ڡ�m�|`���?�����'��޼p��e8�;��I��S��Ȥ2ӔPY� �ՠ�h�(VS�U|�l��̌���޶�f�=����	���q�ӊ�1�qv���4��6f&����zbf��|	9�e]�D���=���\I�.��{��0\l��e'P����S������޾����o���32�q]p���o�� n/�\|y�z�`fb (�����4�t��(��({�@;|h;���`�{V���Z�����1ʼs�~�{{�a��?~��B�b茅�D��D�s��kX|pV��u�m#+ʨ+�-:���'&�������۱#��������^�t͂b�ni^Юn��'��ǌ�U&w�=h�<�,��/;�.] ����̔O�8C�?�C;޸�a�N�H�6�����<���<v��ľ}K(�����Wھ��qg�-Ktduܖ�%U��2�ٳ�Q���=Bq>fP�=dp!@��go;#�i5c.�/v.��:��=�� ��,��W�_��W�\�h�G���3�YA>�*�0`ڷ��ݻ7�vفe�BQg9�b��b�g�x�h���3�gӎ/�!�vЄwv�/7}�h�I�7�@��n����W�}��o� d��,f�}{�}_n��=,2hs_Z����Ơ��;8gR����?2��&d�EdDy�:���<DGGH�����1	"�I��W~oў�q��!�z�2������^� ��,
�{ �^��ǏV�dف�ӧ��UW(��ЌP��<���ia ��g��^F'�����٣	3H���p�Ed�P;D�t�k�-0��)�l�9r����ch~�X~? Tw8r�&8wW�m9�� ���e����ͯn���C���?$n����O>��ݺw�?o�Nj�Nig�C_�C��[�ɷO�^�E�9D:)%'ѝ�O�C@d!/aZ���������O��C��y�nZ��{��q[D&ݒ��o}������c�O���ﴟt�}��?�^��:38n���v���fx�1��:fn�r1>�&������qK��8k�!��փ.�i�ȍ<G�ɤ	^J]�bIX�3���	g�4NZl����0cGG�OE_�[e� l]v��A@�����7^?�>>�U���e��q�F�x�b��e�Oܟ=s�}�ߠO�\�'��.�k6�^�|����M�P�9}�}�����8�F}y9���+Dk���ڕ�7��+�ڕ+W��;�Cʦ۝j�P~P�W��������Z+N�: �i	��&��֮߸���n-��T%aSI�1���ո6�T0��6�4G�tJ'nO#$jGڿʌ��N㶨��Ԍ{l��g����Č8_f�#�_a&i�$����A��Z��6��bܘ_BN��L�mA}����������vY��i�3F��[kB��̙�#_�ׯ�m?������'�nk6r/Ϝ�Z�wIb���S�_�A�i�OngϞl'O��`�O����>�����F�X�сnh0O[>j��?Ƚ%��ݿO'�H0��2���4��ѕi����2Ʊ!�-n�����P44nA9�i���ډ�Gۉ���cG���Q:Ӄ��l����Z��ǵ��X��]]�t;@�x���v���Xϛ���	��8��u�\	�_un���η\ʀ�J�%�M@t�-�!8�v��y[jǎl����>#`Qqfə4
L �Plf���r���v���v�ֽv�o݁n@��חǲ��nT�$m���YŨ����L��\Rv��l+����C�����8�� ����ߟ�}g�L��+���u�����t�������* _�nq6w����r���Dg@�v��?���3����B�@P��ڙC�~x/��
f�b�� ;v8�"���n��yi��̒ "@ݿ;�8|�r���=xĀy���~;�nۘ�\F�8莖��$��.�7�0 ��z C{�v���}���(rB{T�lf%9��3��,H�,��'���O2 ��\�CV��=a@J�Asڒ��^g�L�u����Ɏ>���oV6�V?���@uж�4�L,G�� ގ?�A�>9���Eڔ��1��+���=:v�-�:4�?V(Y�9�[ |K@m�Kp�p������i��v��{�'?����_�]���w�log�۷�:۾��[�4����Yv�����f	=��|M?����V����x�4�����]�~�r�]�x�ݸq�r��?s�t������ڎ�<��p����������*�{�[�ümV����o���f6�Q0� ���3�.b���WFX� $�	Ȭ��O�l�'"~��M��9�_�`;��-?���f)�g��3+<	S�+��&e��B�mj_"��C�7�z����[���ӧ��MI��7T���K/�c���?��۽�w�2s�����o33�������B� ��_�z�:�( ����g�?���z.�����@�1��8�����.�k׮����	���_bf1H�"z�:�Vm�nܒ�?����y��i�.��t:̳^#�^c�SY=��l�?+�4����P*zFz��s{��L��W�i�������b�N򙴀a��;�?�6�_��;m�e��NM�af�v>�5�[G�9��v�:wj��GC�5=|������3��%֎%���ڤ��?D�<F�9�exgnn�@.|~����>�������m~7q�v���k�Y�u�}���7ε�4����Q�m{�,��[ț�n�.��\F_�!;�x� `�p���,�8���ͥ�ڌ�,`�&RKL������r)Slq�@�3�����ݵ�(@<~� ���e_;�^�#=EGzX���,��.��(�Q��th��9xp�oo�.u�o}��euylAD�B�#�ݫx�Z1��8�}+p0߽`{`�" �@{×_�<���:�3��cG����H�w`���u�q%3�Π��� |���r/���. A�j�.
�R�S��B�ub��aU�x��a��('�i��;ݯ����7_99�N�8@w`q�1��^K�2�l��<GN������*;ҭ-��0�ү+ciL �z2�����[��S�>j3���q��e�f�&m瑑7�<��y�<�u ���sg���(����Ä�Fi=B���X����^��˜e�F��MW��bI:a˔~B�#�����|�Q�cp���Ү ۓ'��N?�����o�����5=� �A�r�zH��@�eYY���	�x8[?��Uh.P ��ĥ\�K�i_�t�9.���uy��m��ZuȻ�+�_{�t;�F�����:Sv�������~��U ���D�jhp��w��*#�r����g��� �+�/3��Xˬ������{o�c7�z�6w�:Wf�u��L��;���Z�?�v�HZ���Wv��=d^b������l6���<?C<��������}��7I{�f�A�C ����F"�[>˜Y۪�gRW1��_i��1~O���_~����b�~�y���_�V���؄����W���
�g������V~lz2	I��O�d''�1�<-j�`F{�{u3��6�޻�w�e��?�U�����n�+�.� J���֫����<�[�����_˶�;��kWo �/S��p$���(ȯ�ny8q�}���Mn޸ {�΃L�lm:1 ����/\��׳Е�lu*���v�ѝZﱃ��F�Ͳ�'�"����X�[*��4%(�P11#��y�m7#�П�$Sf�Ӽ�wjLo�n^ϙ h{�rG�-��̔���VZ��ٙ���F�Ik{���'&9�˺����$|��u7�{��i�1Ǥ��j��4֓^���~�GX4��F*�=~�P;%�EQ���#��n/\���$ݳ��������\�vo;w�D �[tB�]*wfȳ#}#�/	�q���2���@�����}��E�A���ٳ�Z��Y��OukT_�v��`U������GA�/��Y�|��`�m�Ϟj�OkG� �93$BS1��|�Wv;j�1�	[.g���d;{'`�|�n��}C�ގ��R���(ʲqT>w�9�Z�&`yN^��r~���j�zC@N����MK�L�ɡ�r_���^K��z�P^i]Q��3������_�y]� �}^�"��7�������H�߻8���< �5C���c (@�K�.���ahE&��*�3����Z�\ƫ%J��Ex�e�Z�����v��Z���Ɂ'�a>c�Ú��N˙�En�q $�o z�`!�9 ?
�po���{��4�ci^�k;�[j��!�]��Kő��IϞ8�a�¿���p-Z�)�������) Z⯿~��a�z2+�V�l�Y�Y��z�^!���g�l�ٷ��I	^J�{Zm��r�8a����'��Y����,�9��g ��,ο@��C����d����S��#�ȃ���F�
�+���e�R+Kꝲy	=�I"�]�P���:�m�����C��S�:�]ZA�9���������Zx��5�{�-v�^������~x�~H{�c0_tFܫ�����#���VJζ9����v���lK�����*���	n3w�>j׮��JA�-u��h�ٶh��AT���b�T�����q�=��r�������̌�:�?�����WW�KBi���.k���U�8��1y��͡7��F�d�5@Z��N�f{[�5fn�k��0��?x���C�k.]��>�����'��{ȍro]>t(��� �ZF>��.�ݼy�]�~�Aɍ`D��{��	��ٖ%�9�@�P[��?���v��KĻ�A͆�X����V���H�'YAr��J��,���*[�*~���u�u�?���nnם��sh�h*�\u7�⯐bz�k�o�J�% �L����ʝ1��;��W,��X��+���l�t�ɣ��$���;�5�k��j��gx�I��䫙��󤾃��E����L�*�f"���f[�=�$���<�����3<p'��䈳���v��)��j�+w��'$G�`��v� \�,�7P��}������}�cW���v��hک;>i�t�.�q�N6@����m�!9⬗�Hc�<�]
rȭ$M��h���/_ �d�����Nr�r<`��g褎1���ZgY�m��� zyJ�9�oko���|)�C^��'��$�����o`��>�H���s��l�a(k݀k�G� q�y �^�!�����r����h����:��A�*4T6��ۻ�X\�� a�x��53W�h���ӂ��'�5�*3&n���5e��&��w�ބ�$�ہ�	�v6�� g��bx��Vg(T�.�m:0�^���m	 ��.���ډ�[gƃ~An�N�-{;����������AL��g��E'�Ԏ;`�:r"���}�F83�<<wf>�/�\Ϟi��v��(n 2XM����c;��J@_�uiL���Yj!y�Lm���]�h�K�r��Y�6�y�<�}p�|t�;��F6W�����~�p-to��-���V!��9��\x��Z�s@�|���!%�Z���S���χ�)��@1 ����{o���y= ��g;����4��;0�d�+�Y�&��%н{����v{��Nh�h�g��w��Vp{Й[����%�ݿ��]�v�]��b�=�-���H�0=B,/zR0Ӭ#��B��4����pٴ�3X�Mݢ�Rnl��@��`�pnr���k�2{�Iʒ3�n�x��*�ĝ����!X×�ϥ��(!�~�v�}�S���&_�&!z�ɬ+�����rÛZ�*k{���x����
c��%?E�gJW��K�;�Z�#�0W]���jʃt�^�9W���]�e��/^�:=ʀݙ[��2n?��O~��I���?k�o�
�ζ=z���ОxR�+$�YX���6u{�����xM�����'�'����0�:�Y�kWn������?�E�x�����c>{V��{n}9�4�ꒁB7�j�I%��_�����s������pQ�S�Q=1M	������d�~��������γ����q_i�q�`�7M?�W�̗e�Ϳ߼�/�E��7��re�/53��ɑD�w��^>����+�өz�H�O^eB�+�Lw<�I���ALnV�f^�
U@��������> �޼�E��{���H�x������v���,��=�ڙ,�ى��U�s�AЧb�rq_!�A�c������΀8�;�>��E.���/���� ����2��\��3q����);�7�m�~���U�i��[3��n�CJI����m��p �ܛ�,Ht��z@��׋���AК�bm���<� h�.��S �qfI@�l�?�vf(�eS�ԎND;9�?go����\�},��E7���t�̠�v�aO��H��S�V�<�:k�h؝�^g�����:<?z�`I����V@�t�a�����cv��2[$�V���k���X��7�%�b�4��&l�""�:_�\��� ��w����?�=~��֎8�d �v��t�vΤ��*�%\N*����-@LG�,X�MgY���QO�
\�/�5ʉ��N7]lڌy�~}Q���}K�M|�ܩ�wf��׼oO�F#��y�*�����)� ��2!?ʿ����q۳��r"��ذT�+˚��l���>O(�����`�{�����̌�+@g�oG��'o�����<�X묑���ʵu(Oj�ܙh�e����e�|;��sg!\pK}���Ix����>���n^��.^���޽K[XC(G�B�m�ǂQ�v�ʮ�ߒ�6uF� 0�6S|�O~cSx�^��`�K*<�-7o�i��^�pvϭ�����Ҹ�֥�;�d&���G�A���LV:��<�⠱��;SgЗ:{�Q�o\�޶=$U��m@u�+{D�o��Ҷ�w��Q�k��>M7 Q��y���Qu�]��@�e�V��S�.w��4��˂k�"��ڔ��e$�2��vm�j0�֣��~3�{ >z���g?k�~�q���ӧ5�
 ={�,�.5?�"���.9|���д��ͭl�:ÿ��=�����Q��q��2�_7�/ ��/]��ņ�z��+���>�5~�(_^�;*�����we�_�TH�ܿ�������G� �h\��p������|�\���4�V�ⓘv&�� �ega̟ac��{Y�����O�i��f��HHw��I��*ʝ~;��i53����?)�$]lW>�pژ>�W�q15��l��f��/�/3M��,�)�����R�:m��Tn�,�=}��>s
E�\3�7�K��f���\��2q����}�g��og��eZgl����i����F�L���t�f9`���;;�gt
΂)�*$����v��_��}�\�E'��Y�(�ɒh/W)-Ӱ�(�䳅|���'O hى��^lU�6�1�gRY����@Γ�õ/��gi�%ѥ,1g�&�4�����I	s��?�msO��m��&�+�V`	��E�>p{�3D�Nooj�{�@˩v��{��6g3�� rt��;��s��j�Ŝ����k�k��q6NŸe��.�
ȩʔϯf��n�t�
_^���3�m��V�/�O�2� �s�}�3��v!�����"!ά�3��i�UV�B}�O&-�#?�@6����&ȥ.�|(c���G^�a�3���:W��R�tF2�pY�P_�;v�@@��+8�錧3n��V;��
f���׭�� їI\��TH��'nM���BcVI�'�Sfɇ��5-�r-HE�2�t�����v�c��%DrF�Ng���&�wœ�s.�#��)�ԊN�#(�S����x��mח�\M<�G;��˱�7����7Ћ,��_5Z �.ι��e@o�K����������x���΂{r�
C���k�����A�&_P��=�b�r���������%r�̭��<u$K���G�����ە�W ����N^s������w�8ʌ��c�^���Һ����|���v�=K? ���:�Mі,��[������������Y�p��	���ܖ�oz�i�����me�v�j��(���� ���/��&�+����]�:�Ql��e���� _(v�/5�My�	��fW
6�][%~?��6c�V'�O�5��[y*`��F��QO���%�����SZg��Q�L�X3iO�v֨���H;�����=ޯ�q�;v$ �ɣG���˗��۷��cGsd�k����훷�Wo��W�e�c�~O�}ȓ{�2�;B�"�����:0>x�PV#<�����;�y���p�G=�v��� rr�ő�o�>�����@t�}C�D�9��:����>�
��_Vn���ٲ
��?�&l03i��&��Uq�N�N��X�q�Ӧr�;�g�wڝ�^�LbFca��V�_bgM�㕶�/D��R�z=.s1kv�7̗x�����1۞�~�v\�Bw��T 5�7)�2��p��^&�1v�ϙH�P-)��]�t��J�Q����B��Q5Dc
��-��
��Z�����*ze���3JF�N�Np�t9�Xۏ���Ӹ��p5��aFdڶS
I%�٥�݀ۥ�t�Q+`ٻ�^�EXhq/��S��v x
s�}�XϗT�:#1�`'n[�#���>��9����#���QT�$�a�h�)/u�Y �}_�3��s�4�ǎ��o
��P��[`h��n��) �a7�G!ٹ��+���>�<M��L�/�9�岭{��g
��R����%:H�D���t>M�
���V�η�y�XV����,h	��� P~��C 9ׂs;eA��*��нEGh^֩��ǎ�~��'��Y�T첣��K�%'C�F�[�T;xehR�}	񰳶�����Z�y�������� �[��s0$�s�e}����֩�hg�_RS��Sǩϓ��IO28�w�v@'�P�C�e}�5��j;����N�/I���A_ڣM֋���}�ȩD���l-r�Y�y��n>\� ��+��&��'�=ȍ/*�;}"gy��C7�e�����4�G�4�J%g�Z�ޙ~^6\0�����6}�\ �G)`I��
 �-�q�m4k_0��g��_~L�e� �d���ξ���6��R���>V=f�:����i�։i����0��6HZ�PK�� ^�����9g��peLP�β�t��U�:ρl,t�_@�����>M�К�U��mb��X�~Ua����4��_��O���ۏ�_��w�׾�^����߾������̙� ޽��:�F�X?� �n��o�=g�k��V~	�O9��|{����W�Zy|��>H��v���u�6�L[Gn�r�Bʐ��Z���6�#y�'�4��i��f��v*�oSUx"?����]�Ν����������;���0;t�pNP{��t�G�_��%m��9]��w������' �ՙ���Q����FY�L0���R�5T�����@���[Ѫ!z:QnOB��/�Bi�8*F-D�A��.��A�S3�T�g�*��~�ɟ����g���6����:k	��x�NʋWXMҹ��k�M�,�Y�-������^�xO�=��v����SS	����ᓿ�%(���|���Y>܀��e:σ .�C���c��5r�A���I
�"�i<��q�����P�;��=r����S	Pb6j���.�2V�
ʜi���'J?���w8Vpag�Ks��D}�F���}{<��R��S6:G�u,�uɯfk�(lgm]�-pm�e'�r��:;���S�����/R�t�2��~*��Zڽ�9-�4�C�0�o�N��� �����GIƾ2_B�e��C�8R�k�2�����ݻ���3�.� ��|���X�M%<�_��C�U��qz��Y��>�Q_��ղO�:4y(��� ����X��X�\g�S�ψ���-z����!Һ�x�q�ו��*�%w5�/����sD�c���Ϡ<{�T^Y<	�\rvv�<8��ҷ֗�b�	��έ���P~��ҁ�Q���z��g��Du�3�Ć�0i�����Fl�+�l�����G������V / �೷SAzfi�u��A�{����r��@������RN������S2Rd����[��V�v�K��.�ȝ��.��=��}�Mf�y*�謷�q�W�K����	kf�w��<_��
r=�y)�;��@;�=M��=�#�ҍ�U�{&�p�^,(�h۞2VMܧ��/�=��U�}����A��R⁽ꢕ��e�:r��q�\���h*3��2��6�˓�v� ^©'�T���w��v[�m{ܟռ�|���o~�~�����w�޾�[�l���_o����h��0�g0HEv=�����k~�^{���NmO�����_	���?:��ۤ����v��w������F��w���0g�:���b�i˽�N��:�i���j�&2y�=���OW�`K�zE�8hw�D�u"Dٰ?~�$3�����_|�~�ӟ������ҕK���Gщ��?~�!�����wj��z�k��"�D�z�-u�-�9���0�����o�PvR�R<�62=9�K��ц7��-�c+A1.�����*�6R��L��$-��V��$��3{�f<�i{��j�������4�}��/�#�X����$\5֩�y�-܈�/&a�`��og�ٖ�;����1�N���ee�L���X#�H�U�=��B����>��(��X|�ڏ3���^:'�}�Ea:�ಡ��(�r�i)�U=Ո�ׄ��Хe:0�QΣu�r�����H]z�mi_B�3%�M��ڴb�b�,K �V�
�T�g��j9k �.��8�=8�Ѹ\kc'Fb��v�sЋ>+�ʗ�HC��,�p�%�q�׎jЕ΅�$�S���*�
Ĳ����#���>��Sޕ"6^�eQ��l���e�b���F����m��c<��رC��#�T<�ș�l��*�"c�L:F��%C�]_��RA�/h�4�][�N�o��lO�/�	ؑu.���n��v�~EL�l��l���р��a����F_�)ܜԑ{��ܢ8��L��q� ��R��������g[���s�{:޵��U��� ��{���t��Y<��ʷ�=���l/��˛ًE�m����d� Ҏ�7��)s~��c��M�� ��	Bs��)G������Lyfͱ��	�)�rB�r��l��̑r�G�%�L{prO���æ��+;��ܴ}e��[�@v���4^
�~����ٮ}O30�Fu��G	k�X�]�;�tF�6���r�a���p;{;�����m�!mtZ�ʶU˅t��e�ʨu��{?��֬լ�F�W_F�k�W�qU+�!�N�I�4*�9h�O��+�[4�����e����;��ɫ�4��6i���3���n�x͓ht�:�jٱ���ײ-�#�Μ9ю��u;��o����<�eu�{hU�zB����7�	=��)?�̇<|��<�(�F~m��	g��ā���Y��7�;�'�����s��'z}�b�W4���=n�8 ��o�,ٚ���c������K�g��.]��n߽ó�m�+1���kg(���8'H���L  ׋��2zp�}���v��	,�}��
z�85�P}�D�w�mbyf����c�j}�%(\B�d���%���kEs�t3���������5��F&��1>�5�n��F*!���Omŭ�Ug��z>2�ٸ*���-�W�#���w���vw���΃
?�p���x����_~&o��⋶�������kc&q�Řn�,M�N\l�P(~AY�^��D�W @g��uܗ@��uOnްv�k�%m��2���"�˺Θ�
��4��W�߶�\  С��y���@��.M��
P !hHC���z�����E/g�ݎ@G$�u��Х/g��./Q&:Q�T�쬳�@p	(ˣ�J����y
���[����/eFڔ��V��UaX'Z~f��|�7�2�T闚�5�'mTt�V�a��M`�wQ�X�M��	������ֶ�K�Z:'��qQ =��1;�dH#v"1��Al��}�t�,��|&/��S��2����X,��f��,� �����Ő���-q��T�Ei��$:C�lY�l��/�-1n���l�jY�-��h�:��=����m��'km�)���ou:�\��{c��l���O��~6���[pц\mȶ*ܗ|��ݛ��H3 g|�Am�;�ڒ�Z<S4l��� ��s�.��Fw�چ^X�6���	lm|0�E�%~�ir���8��i�Ѧ^"���!�m"�j���.�2�XeE%���Q��/��X��8kw����@9�NY��P���yZ���������2����݂b��6`9,�2�|D&����90W79@��X���@e��*��L�Mtb�j,œ����4z��m5`v/r� �<���ޏ�x\ْ����P�ן�֓�O=˷�s*�PG��(wae�{d��1��`rO��\��޷X@��fS�/�<���V]2&$J��J���n9�-e�j�l�� �2(�u��������}�����v�4�4���-ʂ�wP���X;O��+��0��:��)�lf�t�A�9@��S}�6�N�M[����˞�s�<K��{˯����eڧ���<��=�ǎ�l�O�\�����6���1�����G�о��-�v���v��v�{��5@�_���j��R�*�Уn+�<@�9t�A����e=~�x;㋻o�o��N{^����'W9}	��g�Ά�MN�|����U���(�/��o1І���ʤޠ
ؖ��_?k�I� 	����0���/���6���N����k������2���睖i؊�F���W�&�ݍ�8Ӳu3>��M����c3�zv:R���0�ˆ�m&5:.v>.�*?��+3��n'��ۮ�K�pSVX/���
�-_9
�pPfz����ᩤU�Q�1�(.TZ���@L�|(=����En�;� O\;��퍎��f�%ᚽ�y� �u}�a���@� �"��׼�-y�#g&�e�!�/��CZ���*�_�X��m�`�Iϥ����t��h�Iy6f�w��7�]R�ov���:g�#�S�:�+鮐����O��24���Z�C�
��f]���=��3�V������ҷ�8*'Yj%M��8\JwP ��˼�׹�(�6�)^;�[K����v��Cǵ���s�.k/S��ZP@P�uǟ A�Z�|�*�g�Ǡ�P*������X<B`"��x�sm��:��-�ú�C���`�ˊ��O�ҳ����4�W�X+�{�S��������%�r$&�ڼTh���֖_���Z������Ƣ�(��--��5~��j���*7�%���MF��u�`v�r���q�㮭>���O�Q��"������|!?䧼�R��C��wl�9��L[%�zCy̹Ô��.�������r;	���П2��O�rѕM�+2!��\NW��tS���y�����8��@�z8y+[�v���ц���Vb(�V��G��S�	]q�`RP�n���'n�p䀮/ی[z܊�Y���'Oۍk7�g�|���]�
p{�8��U_��]
W����c�ã�����*��$���j��b�_��|�R���Oۅ�?k�n�HxW3�Ǚ[?Z�l��׶�Q�Q�nan��!�X[J���w�T������.nҶ��S�����>�����~�������c�Ŷ���=]�h���V|7�H�a=���&��2D�r�V|hw�8�O�1�JtP����x띷ڇ_��}�k_m_��Wۇ��~{�w� [�5�[j��RѶ��e��r����[2Ɩ��(��P�I�g1K���b��M@@Q�[~��������$"�0B2�6B?cǈ}j�!�w2)�+����h��c��ޛ�v�Y[�F��k(M�Jטlb�3���M��=�V3�'vJ�f�m�zj�aRW��u����2���It�C'嬲v;uؘ�g�z�?��x�x{���&1��L�Z��@B�$�Ȓ$����&,3�JO!v����k_�K��e�q&�%j�D���c� Vٝi�$g�,o���F ���2�z����##M�V�-�7�/K�О:P���׭���H���~5�\�&W�L�;!g�3��i��n"��� <��JBz��N'N�A<����K��գ=�Vi����N%-r�+�t��I���aj6��ףq�S�ò�S�g7��3��<ȫ��w�(cK_���ì4&:�5�V|I=���a8i�})��~�8@�������X5�@r�@²����Pg��*`���`a�K���4��c˷���; �a�U�0�� �Aʊ@�P��7���&O �:�Mm�lm��)�.�
\����t�Yּ�(P�~�\ C1�7-�kE#�c��p�����/����Q��ӄW��z�P^Y.�����͋I��u�O6�(v�-'�.�:뜭~l;�f��h�m`�c�(�����.1��o�/��EG�5�,��lh�a�%|N�^�G�/�up�Ud6/q*g���D������T�J�9��T&X��-�.~��g�\&��O��tk����ʂ���<�C9�s�2\Jۣ.�5�L��?t�2���tݗ��5\*+u���b��6���!e�5����ß�ʴ��=�[��������������������៴?��?j��~��_�۷�|�r�sxb�#ʮq˽�r%@]g[��5�km��Z��u�+�'?�y��?�����'��~�ӟ�s׆�(.gm���z_?�A����ɰ׀�ݑY�@P|w��c������O��2`���������ھ��a��W��N�<It?���ݾ��=|�v�T�w�}�}�[�h�������w�7��M��k'N��M���t�u�N��޾}���o4OSx����o��o������������?�'�������}����k� ����l�f�j[u���Lʨ��wY�Uޣs��X�H�R��zX�L��w22�G�E�@!�鰒QuX�?��obz�r�Q�Ms7ё8$C<�� [;��һ������d4~`b:<�Z���N3���7I��>��27=����Z�I��R�*�n�7���ʤ��9��x�\7�������
��v�í4G�M�+��G3a'�_��m���\L,?�a�s�{:�/���{���Y�Q��2�"�Tv�r@�f�A�Q����ڸF�V�U�\v��H�����&��TY�}�� �$G�ďd@C�&��!(K��n�l�(t"i�-�������c�����Y��yfV�:�k�緂i��܍4&u4,a;���M|��@�I�2��$􅟕�����IZ�1���|��0��5��� >Qϵ�l�ZV�Kw�U:l��#=y�lF�J�QC�|N�a�ת[bॕ�����n���t��]e��[�N�)�<*�8�k��x�Fp ����5��[��7��;�X�
�Oy�,e�E�?�:y鲹�ϬgUe���V��i�^Lt(:�Uv�s�9�!_mѓj���
���0Zc�F��; y��ةBV;^���?%4����J����0&~2�XAU��i�ӭmm@���ɞ%0*`�A̦�嚲��u���n��ݤ��؀Zmq'�����F�RvlG�����I���qx�U���u�����!�|�~�Sk+��T@:�0�l���qN�S�$�Ns�8�Q��
k�u�-w�����k�W�<f�!�)c]����0y��.i�V̺v�k.������ܾ}�}����c �������~�~���O�q����Pƃ{�ړGO�X�o����=i�S�]�l� [�x��Ӌ��~��g���+9fK�i�uz�+��U?�uRmV��f�T���0��k���V�6 ��v�{�=}����;�Ξ���7 �E��ÇǄ�ݮ]����y��^��A���!�w��o��N�>�>XnOV�I�v�p�j�t�Z���
7��s+�gϾv��k�������{��������m�5mC�9Sݖ��DFf�À�7�����'�&�4���û0�(�X6��q�D����ĩ���ƀ���W3r(zB
�§-�`��.u�T�^FKڱP�u��l�L��(�%�ʉ[���3�����6`2�Yfky&gTy���6
@�a}K��ׄ�
%�ً�y��Z�������^��;�TBڑ���⇕�N�Ί�3�t��1���tziPN��%�4#��̓�Aӌ�	��ì-�L0���=����ގpj��|+�aq[6
4UC���ϼS���\i�V⻄�����B	��>�%�BA���,mf��������Ҏ����Ӏ��I��q;s��/��;���oo�d^p�:�T,�9����Pl���Mz./�������Dfc�����nnb��v?�5ڹiΰ�����#b�\��0�fGL�ҐsF3l����L�6c*�>�~��k۟��$d�i�ics&��t�i+��V#�	*��S�l�*�s�ƽ3���挡�"�G�C)���\���9Q����UI��D$9�NY:�!�㲝Q]U���K�z?��'��������ʃ�����+X��kQ�8�:�����7-ߥk٫�K�#��Q"�'4G�w`����M�~5y��nM�A�=�JGQn5�y�D:�x�i�&�����	e�8�xɥr��V��ʇ��)K��I��uh3?����6����������}��)<���T�D�������Fy� ����h�k���m��-M�ve�tk�G���R���:f��'���4�1@��@e0���@�����w��3jS��Z����+/u��W�����:��۽_q�V*���ѡ���>�:�$_U��~C�\)��� \J�#�)k�|r�`��#´m�X���� �|�7Xüɵ~ʐr�I���I�n+X�M���|���'�~������|�?\o�n?j�.�j>��>�ŕ��|���������U�ُ?i�/^�3�ܼ���z�=X���WX�걱���g�޺�>��ǀ��~�'���W�k<H|��v�� ly!<��#��.�j��ڰ,uٱ�m��|���C9S��n��v�.���s_�Ю]����B�o�'4�i�=��o?������>��Z�q�^{��i{��I�L�\�9~�Hfy����/_o?��?����G}N>W����ڍ��ڃ���6����[��͏�~�@�Z{x�Xq#mҺ�D�J�W]��21���R��טHm��{�A�/�S?#(0(=���P������x6&��M��<1ɴl����4���uT�˄������Ҧ��fY�h�s��\��n�W��fM��_�k~��-�-���%���F7c�\�]�b�gF]����4V-e�WQ懻�ZT�=�I/ ?{R��U�m��b���l��\�p&����Z���"���y�(����7�� �PS�_�4��ĳ��q(�ͳN:���y�_�q���N�Fc=��k� �Ӡ��";S*��K��l���ĥ��'=:V�HU0�|�T�S�*�.�k�ꡬ��m�y�Eb/�H�·�ٳG�����j6;AǄ�.z�&]lfJF7h��*�*�t0<���ӳ-xf�U&y�S�&���o��3���[2ߧ���3d���H:C��U�U������#i��'m�k?%�5?�����X�W �M6��Z�?�O��,��uf��_�%�Ɲ\'����I���_�6�Q�[�4���<#��r`0IXW��3�(s���l��X�"-�九z��S��k��0t�̧��ʙ/��1�^d��x8��-�YH)����F~��4���1q�*�����T��G?�4m�� $@ۿe%��U�HJzv�-��m-��f�3ߐ��zt�����.�:�[Aw�^,�M{���z�����0
�����~��K��#�g�D^m�>L���M�<`�9�"��-��KH�ͪJ����Z2�6�5)^�̻��M7�E�7�yP�����Oڨע�b���V�c]���x����Ŏ3�7\3�ڮ3CN~U�(�E���?�d��� ���!������ ����?�л���y���}��zgp���Q75"����>~�8[�\�J�[�0�_Z<t�c϶�'Ne��u�v?j�ٲ�b�v1!tX�낒`��պ5�xoG�\�C����|�֙cA���g��^����~�K��_\l/\����������H�����u��i���k�n���R����c/|~��n%�=�䖎K�����?o׶�r�Zh��u~��QNzq<b���(r5�a1U���.��\bfE�������"9S3��[I�v��Q��l�	���_4�o�b~~�Q �l�i[}��=}���>y�֞>n�O���*�V�&��gkO�O�3���ȵ~X��W�u������Ou�N�\�ſ���:��D����u����'h�]��RB�y��Rxu�-�٤,ұ��~[}|���>L��o=[E��b�o�buǽ@���箾�>���K0�m�o��m�Z�n��y�J���^�'JZ%���Uіu��m�3��_j^�\���mr��6�q}��3�rV�#����q{৤���~;mW�=����3�Z;�R�EO�H�� ��&@je�I��.g/z�I\�\�x�%��5�O�Y�H!�Ƚ��'p0��Y���p7T����["�w@^�ײ��x�F��uƎ#��Ya���sΈQ6�O-����í�K�R�
q��W��0�Q9{#��ى \����(*`T+.�8/����E?`e��&���^h���=\�-e�X��K�`N�=�S{� qԇ�5��p����o7���X���/����$j�t�1��~��"o	�<3���AehrF��X����F�ȅ��\+_]F��:) &�L��1xʶ��QI* n8*�@������ե�SGc�^v�'T�r�U �����\WYS/rM\��;�X_Xy�>D��:y���7����o��ժ���H�7@���s�-4��R���0���� ��	�=W�x�<�c������Y˪K�O�'O��_XZ�L��v�Ȋt�/oj�_Z�v �5�����/ku&z���M�I?-]/�ᩱ|\��M��E:��l��� ��5\iHOr�Y�yZtk\��4h�%Q=�e�ڮ��F���3���g:;l�����V��U���!��{x�v����R�v����n���Rʉ:c|���I��te�A�|mQ����6�{��E_�Z�::��rf;�x��g���d��u?u�3��|���v��8������r�*a]�vyށ̐uH���Tz(o�r�Ǔ�� ���2�����Δ~��_�����n���������e�˿����8�|�ݹs:�?��O�޾y�}���}�{����/��џ�?��?o�g��������G?n� ��-~���nP�|��ӏ?i?�������������'������>��ݺq3/�yJ���(�v,'�,�(׌�e�����A"+� N^���
o,�*�Q����9�?w	95�ܺ�yU8B���ׁڞ-��^8� �u 8y��� �ϱ[k�/���z��j{`|������z�k���%|�{ZaM�g`n�;PT��P(�@0C�q�{���w�y$I�<�I�Lk��*�O>�<OH�<�]{�u�/�U>m���ڣ��.�)�F�6)Ӗ^
��9V���md�N92�b/J�깗/���~h��l����J�����"gț.��J��
H�S�~��7?���(Xf��l���S�r��#a�(��#l-��2xٵk� �(�(��?y�F�VIy�y�9��Gb��6�V'�27%{m}�=y���$�<�~�TpM����v6y�>�R��O>�X�$_��3]�XP�����)�p�o�j�������y ��*
�ȮgPD>� ��sW2x���������^ձ9:+*��3�O���'v6v&��<�e������JV��r+�D�Q?1��'f7<o�H�%W�b�UTl�1�0������,[-�[��G ��Q\�|��t�s�[i����m�4g|ed2�N'�U֣���z��R\����.���=����t[6������ 	�=��}{O���.I��2�����K��Y���wϱ�@���=͗��I:�9q���+q�a�����Y��$���Ke~Ƚ1���J`��,��`F`o%w�^�&4�?mK�R�6��Ys ����Y�[]'L�>˴�aO;v�gO��\`����]6G=;�1_����+�e,o��E�We5��c�s �L\��
��`��<�։ 3��,�������)pڞ�`[�ߐUv\����k�K�}�^kH:���6�-�-^���	`�� m��1V8�Cfm���B?�٬9'���$�o��ᬷ+�ʨ2m��9�x��3���i_��%L��@��փ��F���au�6�&��>��FM�L�r�<Ì*Wڠa��*����4
�� ���>t��'?o?������Q���O��4?|�A�����<zخ_��>�����8��G?�!�B�_��.���ol��s��'?|Ԯ]����O�~
��~�)y��}`{�=!�� L�meH�)�������o���a��֍.\�ޘ12��5�LŚV*5�mO�8��ڈ���ǚ��|v^�^���܎F�z��`=<i���׌�wÐ]�����5n�?�{�p�ݛ�e��MZ�������g�m�����E��y�����&�k-y\���T���lx�������kS��r���ϙ_@����C��#t�S��e_�9.6Ϻ�R���ğ����>����	B利���u�vVd ����y蠬���9,��f�����eG����_n�J�.?�M�:ox�,f�:��_ ����R1�uO��땽���#Am�a��GJԕV����X��?��y��Ç�x�۷���n��p&Eѐ���4�}F�O�>i7��ow�?���̳�s���(est-���%g�e͠@��Oub���C�6x������1=yT��}Y��ȡ�.,C��7f����P���$�,�������
p�$�T�-@Q� F�1O'g�j��A|�H�����(_�s |	/���dH(q� ���%�v�㲝��w6�|5֓3�1yY'(�,��c>���L���zV3�ʊː�5?�����ܙ:��j�G{��Ec�c��O�+��I�e"�����l��f�P�LB�y�G�-���S��d����r�Iy�Gj=���{��r��r��Aă��iO EG�(�J��e-	�K�+�d����\�����n�rR �O����ړ������C���趡���m	�Z$Q�M�]
Ȃ�8;�*��p��ɓ'��#��I[G�)w���o0D�
z�s��Ƞϱ�E����G���>�Mp��G��o�S4z:��~	��̜�.����Oٷ൳���^An\��s�^� ~������w �� �O�t[��0VI\����@��C?�@��`��ų���_���_Ү��3�)��3 zʐ� ި�l�4 6�돍_=����3�ŶE�m[�Xwg�~��D ���j���Մ�r�홠9j1灿h�`���m��v�����ۯ���y��8y4�e��)��宏��G�XZ�o�og^;�Ξ?ӎ;L;���ݻ�� ���?i����v��t92�<�Eɕ��;����}Xp�Hږ��
��!�o�1��+ʋ[�Uԇ�B��(�����_ ���޾y�����; ��Y�v���@��@�;7o�+�.���}�.Q�+�.N�������^'�v!K~n[��j��{wۭ��ڕ���Y�l����/��仆�5l��^�m�ۤ P��ɩ��¡N,k�8�<�n�a1��ƎG���F;����F`�ǎQZ=�vc���A�����Px����v��J;u�p;{�o|�l籺~��/��-h��}��gOk��%�����i��sgf,�c�m�i�%}�Vb:�|8����9�|�Tl�^�W���͆}5m��Q���	!��0K��u��Ǐ�o'��l��������IW�����5��v���v��J;zH�LZ��K���M��/{p�~e��{���}m�ޅ�o�B�<M�M��/ʻ�B�^1`���6D�o��;��f��f{��eKh�]�J6�U{G�}fn�z<�=���.;�04v�t@��������n�}�V�<\.tU���E� �;w�77�'�3i�3��̭d�y�ǵ��L=ti���v���v�6i�y �p6Ѽ�ʌ3I8����oyIe�B /�
���yu`vf��e۠�|�t�ݾ���D�޹+(u&a��1M��#m�As]l��S�n9k����vp��7�)�n:�,mO|��m��D�N�f�����P����@�*/�.��^�2 ��ܧ /gn-w�9�!4n@�H�}�ֿ���5�G�d��`�m&�5� ��OGc���C��u8�0Y$� �[vyt�<4�l<�n@���'�%u��F��E�iM:q���bU����: p��4�Uuv�z�v������[�N�: Zgk�Q Mo�9i��a�<%oʲgd�
"����ɇ�R������ S@������S�v�v=[<&m׸�e?r/@M�J>��3/u�?��e�����3�gͺ�]?�֩A�K�D2��HA�Y����J���\:8��<$$΢G���%JY�ˤC~	@�v�4a�)[�磧J�8 �^i�Z����ׁ���2���:c�IxM	H/�P�?�~�(uSQ����cOvVS�C��_�	x*R� [s�lԌ��;����M�^�<�M^�w;�t#Y�b��~��L�mkC� �׫l���FQ������|>���O�:�ΜK�'�|�\���w����N�>�Y\?�۾��qm����.����[�X'�:�νv��f{����豣���׮�k�n���\���]����'���[�'��CJ
š�+�w�	�jz������E8��x?fU�W����ն�V�3WS���h���2�Ǻ�A�u���G�c��\�1P��y:a;b���kO�u�h��?�>���&��g���~h�|֙��"�����X+SFL�����y5����������(��SF��j�h-��0A�\��B�����3�k��'Ś��ak4gV~"�z�7iY@���V;  ���B��Ν���Ξ=�<��(���|��̩���ĝ��i�~�ʞ�^�kj��X��|�X;}Ь?���Z�y���v����{Q��ً�����pQ���b՗���Ծ=� ���$`�����R��̥���?~4�	<v�C����i�s�ُ��> ��[��`�����c�����C�(�����=�-�p~=i��oh�u�=�i�r�!�66�I�DQ��%�,�lY]��O}�&�kj"
�tc02�<��>��,�i�s��)��r
P^�z3��Y�����Q��Q,*&�3M�ET�u���3���T�v5;�WySfg�n���{ڮ������>�=�>^һ���og7��O���TLu�"r0��	Vo��������"�V��I2�)_�p�e��d&M;n%����*�w�dWۥ+7�'�^jc�]��Y��� �Y2��I������c�[Mܯ9�g)��A`Ȳ��������!��F�.P3��
��%~@�sw�O~/R�݀�u:���ҥ����`�Q�����>%+;4���i�#�ss���b����~�������^��̀�h�W�%��  ��[���
l=)C����z�"�����͛w3��Tgxkϟ�T鰎�ֻ�	��9�˯�١�5��Չ�xT�3�ұ.��9�}��ٴ��<����� 9��,��-�J�4;s����}�]EV�]���B��E������%ֺ�f� 	�7?��N��:��
�	݂U��8zdX>���de���R��u��;	��ߍ|��85KY����!�נݣ���?3tf@��+}f i�\H�[��vq������=��u��1�Tf��n�p�δʕA� ���=ki�UN�p���w𺺺�@�!r}�]�r�݈���޽{���O�G��ƹ������[k�i���4|�~�ϧ_k5?�z�� �T��@�ki���U��oК 2�k۰ Q�g�6�w +H�]���v�}C�ڵ�Y]q���y�Jw����λo�=��2�^gP}�]�p��֫'[d�o��XI0�)T����Hb�E�c�{���E�������ܗ���&q��cǏ�w�{Z����ڗ�i,���}ɛo��N�<��Xʠ������G�g��D ���\Ovee	=�m���'Og9s���~�x³ȩǒݿ� X��v�'��-u�W�4r�%��:����K�y�w||ε=��\,خH � �w��Yz�I��}�/{���=��S7b���+��_���򪓟�"}R�czx$L^tmb>u�z���N���
e�V���-[�aJ���%���g��t4q���W���3 F:|��r(�'�F��J4&��sK��0�H�JyŌ��X��_�cG��w�:G�=�^?/��o��~JO@(���~:@��ӓ��{��:���a3��{���i~:��`Ý$�C�J��׭e�@A�s�}�@	p7)��li8L��e���y���F�iӧ\6 ��Re�B����g�Nz,��Y���?�̳�GQp���%-�}.ON�̸~��eA�I�3��8|���Jw�%����`K}�GU��8~{��*Mm*��3>,�.�0����(���/`�K�3��u��jf�2
v;�4Bd�U��=q* �H�D�6 �ȳ�*V�h�e��i��Qg�g��X���_+xy�T%}���J��:����lvZ��,�7 2�M�Q	�>~��� Ư#�IL�^%�N��@u Xh3�V������Y������v��v�����g��sF��{Q�hY ��S7��گ���k �Qy빢+B9ؖP�)m穅xS���~�m�)�k��������[%\�����p�z����<z�r����&�H2�������$��(\��+T���,�@� ���*�4�[3d&&�Τ;3I�8��n�7;}��(��?����:P�C�%�[hu��U�Z'z�
���`֎�b�@�t�Z>5�6��.`S�x/o<d)<4;�'�	A�L�L���o��^l]�z�ݼq?{���e��>xÄR;+���,��v�u?dD^���?t� <߃n�X>z��4:� 5%e�2�^eZ��t��Zi0���_��~�N�����;w|Iw=es�}VS`Vx<�X�V��J�V�M���`��)�@�W�u^g )����� �G�I�v���ܶUs�A}H9��P�h����._ǽ���&�"8��N>�:y����Y���Մ� ����i�$�P�S�{�l;pK�Jo�Y��Q��7kM���Z�+�����/La����uu��a��>�� �')�N4���~��	U�ڱe�<�;c���C�)�H���m����<��p�'��Zٳ��e�� ۃ���3��º��=�'�#�|�5���z�]ܽ{/�^�*�o�y�z��(oϨ�G��x�в�@��i�i�ν�/t?y���/���I�� �'x~}�'��vv�ɑ�9v������(�;	���b#� i�;_�CsjS����#n5��W���um�:���*������3\���90�b���}����Z��u�|	�g~�M�o�j����-�?n߬-!�0
�Ck/Kfm���J�S��Ra�G�J�Ul��z3l�ȿ�+=�S������������?ẍ�Q�V�&�0)7Dޞ���
<��3a�HW��*\�%�Y�g�
�3���Μ<Ծ��[�w^�:K{2�R�vJp�=M÷�a��=!h�qgx�� ������- +���l7���!|vB@(<y03�+�������V�屝�T�M�m�g�e۷�X?�^�
�?������3#�̰�@ }�ܙ����T�=[��e�E6��<쿦k�� �|��.6���3(@)z��[g���q��֙��h�G(�B[P�Aa��[o����Mu��U���.�$��Y<��i�o�?]�mfn�&8��rzJ����;v`��:kf�Xp��e��<��;��¨�Q�5��F9���y�Vp�����Upt�9�t��W����ۥ+��'�\�y|���r1D��rF.�m�/�T���`�����T�N� 7gU.��5W�MfP�����x��Z��w���u$Lz�2O��kn�m���nA�O?��}�}�w��X��D8c�S��I��Ү�a�
r^�q�y��N�m�&f�-�of@hp#;��K���t�7o> h�l�}v%���2��8cf~ă�ꡐ:����J6�Cϔ�ϋX1J��r�-u-C�V'P�KɮdH��a�غ}`�#r�9� ��n��^t�l��W��s�܏Hd d^�Х��7Ց��x�7���=v�s�v��/@��;ŀ��om���&\��ngI�u�JM�(:�|U�t����Β�_��ҜA����l}@�	r6f+3�~r��ѣt���;����������v@!�	�]sk�/�������:���lٗ(��t0+@t�v��	@��I����MyL^q��؁�t�w�k����Jg[�Z\�u�pPE��)_�'�_��k�c�p�g���=
�ȯ]�=�JЭ��)�*϶�������G�ϿpXA��_�x�=x�� �}��󧲂��l�]G���l����S������gՊP}V��J�}Ix���w������I���� ����֡Ç���}�����3���v�s��S�9�'O ��akA2ʤr�S�G�?����a�+kXu��m��>�Q���� �=+{szA���ӏ9z�&���`�� �S>:x(�Oo�u�;v���K�L�~�d�샼tI�\D�O��f8H��/?�^�M�F�|$2v��!�~�9�ݍ,���|l���� =/��/yB�3��W��z��[��#�������� `�?fG�@�i0<�N���₶�_����R0��6Nw�K;�u��$~>;zĕ�C��õr�n6����9ΖGis��tI�4��j0u��e&s�O�\'�2�ݫ޺N���z���hc����p�������}b%d#Ve⿝He��G=��yA�DLp����טbA��͗�����~��[�M ����iq��t�Ea������2�у#	�p�[�o�7�_e��g��o|��gv��7��߻eI'n'���K�7qq���Ψ�(E!z��%���G�XX��ƙ iG���K^������L%�ݛQ����X�#�x>��9�l��_���~�a�#Gd{���!�ӌ�O�3j}ܮ]���	Xj���i�h���:ƻk�Q�C�;1����Dq԰�EG�)nU�>��[CI��u���t�9gn�����2�TcI##� ��*�Z�uK�  gU��f#x��Q��<�F��tx���|޺u7{{="�Y����
X��e��NL(�E�&;��g�y�m\���ŌOؚ9�Q/��e���\`� ${����B{Fg�ޟ���v��JZ�;�LZ��:�*C��u�������_��T�=z�Q���o;�ǃ���mR"x+�9�E֘p�u�i�Q��q޹�]���~^�̏'Txd�3Gv���5�6��!d�8U���bȅ�4	t�}�� i0/6<6��q,��N͇��</��][�I`�"�����,5;�����y�qpt�bJ�@�b�jc�R��≳O�q��쏇@gc��4����"�u�zm��?y' ���uis��g��L��k��WX�謴�|l������gq-��\����u�����$ukxLt�u3��d�[cg�� Y~ B"���� n�O���/]I���3I��m(@���]�˳6��G�F��K�Ҽo�{/�7�6�,���D9�^�7��v !���	0�2=����2" �L�Mfn��
'(�ƃ�k�ƍ���K�H[w�+>+�z��.�a����	�2@���=�D�-�n�.y��6���5�s@�m�/�f`�@Γ^�To޾��4�%9=t�}���5��}�})�����{BzԵ����܄.��iRM�^�r[�Գ�V�T�W���2��E���|�޸ڤ���j�9'�\��@�������$��:�0����{�p��;k}'��寓/�{�A���M�L�a����'���~�1�ց��꯲�R�؄3�����1�b��B���-��0f��.V&��㬩��r|�f�>� ���]��3?�>��m��/�V����V�#Y)v{�Q0� V@{D��qD��b��������y8��=�v�O�['��7ۑ�[��)�
�R��G�cR��Y�u.`�R�m��?����ۇ�ɱBm�f�D�R�c*n���ol����o��g�0�v<�C�s�*�E[��2�=��y>�����j"�"}1ģZЁQ�u�ـ��7��^w֪h&�f�ff2�.���Fz��p��w�o���3�T�)��	`��ތ��L� 
HEu�q䳲w9�|�y�[�,��F:c�n�:A-�#���`�5q���5Q3R�Pa�=���\�7 q��R�'Y��f�cT����*��?���f�e���0�:F�9&3��[����tn}��ٺ�+�!3���hT���K, �M��p��0�33��+s�a�Ӕ%�����%:~e�=�v>v��}~���u�^{��'�]�r��Lg�?Z�v���:N �r/�΂:�*�u���xy��gg��@�J�����l�Q�������
�xHg�+/�����k�'��ׂ3`�Eٓ�����,'ޖH�	Bj{A^�1I�J:�U�ngM�L���`'���fV�N�x��+��V�We ��z�N-�oI�`_~�됉�������R�w����T[(�� ȯ��T���l}V���K�
��"�����X��*`˃�KNg�Ѵ��i��]����8��/��e�G�n��x��yx6l��e�6o]�	��#;�q�sa�uԿ��e�^_�~���u�ֽ�t������g;kg��n*�T�pu��3�st�ډ�����T����0�s�pyY�.����<��r9C�sа���:�S��;w ]��>����h^�c@�ά�-M�LW �o�_7�[�
�u��0g��[{����<Ԡ�Օ�������-z�g�e��ۥ�K��g�]ά���Sʂ$�^�X��[���?���E<z��G������J���7����'E��ʹ%Q��AzuK��m�ՆP�-���g5e���A�2��e@t�A�����j�_'X�}[p�oe�
����k�-���"7Оv����ڒ{�a&����Y����p_q3!ß2�2Z>�{���|�k��Ƌ��>z��^��>��bڮ�`�"�d��;��$�"��9�y-�������MUo�wt��@�)q�w5���~�:���>n����=� E�G���8Ay�غ�Ϊܷo�&���"P�|�}&� ���>���|r]@�	<'���=�+g���0{�6J_�VEq�E���q�t�O��E�Y�%h�?D�~���,������-z���en_d�Z=�u��i��@ɺ��U���a��/�j����>fϭ���񈝧�[Gۄ��"?+)��Rǔ0�5��lE�a#����iZ���=���|��7���c :a�{ٜa��{t־�j���ˇ�����}��r� �qF�~q$qƣ��|���{Pq�Y����8
����Ս+��@�K��Y��[G[5�z!P���/F^�5G.���u	}�}D�������������^�G�ed����\�so�<�ڵ���u�>�R��J���Y��wӺ��亳��(�(���n�v��=]���qk��zm��`GU�C�/������!3��S�Ip�w1K<�
�ƞۀ[�fn�?E�#�%=�����^�n:f@��*�%�,�^>�JZ�*l�pn����r��F@��>�<*h�7�ICЀ���2��y�&�C�{�q�d���@��J@`�[3�(J������;)S�3@�g?�e�l�( ���t?lr�ݺ� �|�N���,�+�RYף(i�t���-n�ڝͪ�S�R���Ǻ��E� CZG�v�� ��C:�۷�W}��V����i�����u�� _^�����ݝ�1y�?�$�7���,ϥ�:$���BR���o�C�`����|�Уդ�A�/;^�t53@wƲ��:����P��d�"�_�={A��Yp;f�ܖ�����H��a��y�� =Ō.P��(+)��#��	v �~ug��kn��H������; [?� 0-�;cGg�돪�:��H���(���:|�h\�J��޶]�p����;m[%Z��*��2
���>ۮ{��@�f=&g®]���s���8��vڈ,�f�NS�R�ю*`������CY�s���m��O �e�Zi���`���7�k�WVls���	}��W�MC���ᙬ6��d���v��/4��L��<]��"��~t�"}�#�d|��3 9����gW� ���϶��C�a���)��^Ywv��w <�}�"Wk���'}��z���$|a��[�zP�*@_�t�{��:����?���n�L�)����pmG)C*9e���m�����
M�`)�7o��@�3��u���I*�Ʈ��E����:��Q��[�D��f�]9QK��'�r|�܋,�p6��%W��غ�P�G�*���Tۖ��٤^d�㲿��d�I�|	 uf��`��[*��l��C�βX4�"S�I��~g��o_Vu��$�����
`�d�p&\j�8�c\��`�g>׺O�v��:c�̭��V������n� ހ\��:Y���~3�h=���/ֽu=�<��hg/��� ���O��x��囙��o���^�����E3��N����b(�	�����{�� t�j���&���ϸ�t����'��G�����V�'��wۇ���s�*�p��A��c^x�!��#�J��A�[9�tt�(mT���`;o���A���ls��,�����}��#���O�7��Q��ep/�s��&�>�2��&)av��(\��'	�1z�.�ScAQ��]�<-�o���ѭ
�{�v���n�z�~����/��'��~�O�,n���P� G
�RԄ�ң�&/g�̪xԩ��{=�ɸu����z��F�x�b�ƶ�}�+��o}��ۿ�������w�~�Y��?�~���e/��< �����?���x�^�d��B�o���x�|{���Q�PZ���՜�(�Р�q��Q��=�M���n7pU�6\�s!R��w��v����z��{�X�q�]���k�'m���v�5�_�j��z��(�C���7Q0�M�����AV�Q�O�: �g��p��|���ٟ�M��2�s�nai���dgMz�S��o�Y�+͜/7�ޙ�u:�U�le�K��)%���k�[��_���Y���J00f���JV����<�h�q�~��L�i�Ǐ�'�k���2�=�	��>,��ϝ���d'`l�������ts���ȅ��k���"Δֲ� qt<�Dcq��}����t�o�y;0t��.�oA/�p �D��z�Ly)=�H����4l�9��K�o�~�}�nt�E�טN��KP.�:�(>��x�g%���_�s��Om޻{?Z�"|�r��o��oR!-��}y�Y�zl�7S���{鞿��k�?�������:��v|��PKj8ŗ���(�N8Kٱ��L\��M�M����s��e�~\��E�U���%��vb�������Ln�g-�QA�\:y��z�ͳ�5�ءt����Z
� �Z����M*d�6�ھ �Q�=�����(c/�L�(�YݑU�
����������C?�@ʑv��������{���'�~֞����~�|����o���7����ٗ-�So5�ߑ�L�`=��mFF�J
<�jq��R2� S��]�O臯����W���ꕫ��� ��o~������o��'N�k7���w����xEZs��s�XVY�"t�����u�;M�nS��Mm1 iB�/�������֓ܮh>n�q0����=���nW8��4p<	޸��Y���o�?zH���g����A�-AЦ��5;�������aM�y6��^��~Ҍ�-�֐�5�i?+� �C��sy�����W@�7���)��V
��/�Ϟ5?��/��W��cT���EpˀS�:c0*O�v��_XϏ}�n�ڙ>�#�@S�u-�ri�n�r� �	8�W��Mo����ѥ�{�&����{\������L�`'��P��C��m�m���W�՟O����ـ,U��A�G�Eb��WQ<��K9{��%+���Ȇ�|�J(ަ�� �8��0�������>|�����Wp�h�=y�d�]@)|��?j���ۊ�_�r�����m&�(�J5&�B�k����I������U�]�fC��Bh]N�j\Ҍ!�0�p�-���v�!B!-2�y��N�9r�-��2h�O���N�cY�qn�fb@|��r��3�����/�;j�ȥ�z�����/~�~���0w��q/��s\%q&F:�/��r�Ji#�2Y�*#1C[�p+�ܽc��nϷo~p�[_���Ƿ�$'������9�p�۳�'$���/�l��ឩ�P��.e��=r$K澈��YT*9;_�������r��3)�cYS_*Q��|)�a�Uƫ�U��I,���-x�ϝ}�|��ڲ�	�勍�O�����Hn}���IE��r��
��4.ϭwg9� ���s+ �G�?�83��(8�k����Խ�6�j���_=��)�����W@���	�6cg�@�?K��ש�ţtv��ǳ-ӑ��FQw���b�l�Tr�O<<�0pd���_#��ʬu�M�"y�%�̀Y���nb�o�W�x���kiޅ�_x���8�ΏODV�}�vg�LO]�@p%��>x {���3:��!Op[��_���l�]�u�@�˿�3m~�$����_ ׁ�+�w������:�"�P��>���{�g��,�*@����Y�p5��)?���9� �֏8��j����>�f��H�҇4SA�� /��_�U��e:�������t�f&�eC:�l��d_+�G[��<���yX�R x��I���:�g�;y��N��@L�&����yP:�'w\#;�g�dԶ ��q�.�"��)l�T�o���P�:�H�דU'擦k�9�w�~���oB/�6���"ȑy֓{?�n�n�>���#�B�����>���ң���W�k����7����ס���=�u�W�oi��M�k����k�������+Fʌ��A� F�b�S��~�팟}~#:�o��{���k��~p����no>n?���w���-�U��u��[��J��ޤ��'}s����o����^�LZZ«���d�>�B�SV�3y�_��[Z쳩�-��6��Q����VבM?@R��j��K}G9�G��G��z�p�uț~�����Y�U��j�Ǉ�� �� �C�-�]hxF�l-gܲ9�{���cW��>��kd\���[&��w>�C����'f=}� �2=.&u��Ǖu1���eG��mҭ��*hN�+�O���j{����*�i�i7n�k�i3y!S���ҒG�}�u�UR�~k�򼠍"'�����n?����  @߿}oA��A����� �Z��_���q�#l	�*}F&\�x�D"-A�?�����]x�N?ؾ��w�?�����|��~�~w�}o�}�����7�g?�8J͎:{K�����T-L2=
7��/�na�/e���3�ҭ����b�R
�K�vA9X�g�`K��y8q���q��D���^�R ��r PQ�IW�cY�'�qc���w�W.�<��V<��K����|�����?ho�����hJ��+W��Oڟ�����g���Ip�Q0��Җ#D��K��	EM�-�T���	̛�uU~����86�bi�t���W�
��̭�v_����?����6p;�=e��/g@�̢o�#��T6�����7�x��=s&�e��Pj���� �%B�\ݢ#rO�{�����hQ%o�o�����^�.w)���rvso������׍<c��KO{��(_�eI�Y奿��j�k�_to�[`<5aum5�����uF�.�w�B����PƗ�[/^�Ll����l��,��W,�
:��]Zi�A���FǱ�=Ҏ>����=��po��W欭_����H�G�y��C@�{��e�m�#w�-3�����J��A1�G����g<ʅr�<�����E@��@���|a��{�}q�d�.?X9�6���v�G�:��vu�Q�^��)���N=`������D�l"�0�H��9�,���i$��4�����isȼ{� `�O�����
��g�A�����+Ξ��R9qj�Ǔ+�ȥy���I�^^��N,O���Vh���;����*��}s��'\��R[-<�ۗb�ʽ2B �]3��a���mh��~�D~S.uP:����K�W���C@#�Ex�Q?ʷz�R�w�_�,�=Z���%t��O��z��J)��wY_JԘ���Mg�D�"��m �y�n���`zjuUF{ߓ�ۯ�]��o�~������}�����]�t9�~�Ϝj������}�����#��3�a@�6���r@o=�ժ'qn)7�P�`�ԉ�A�@痴�B�@��C�|�y��~�O��3u�'�n�3�����	��ϲ5J�DF9J����D�ȯ��\�?�Ms�t�{�O�l�;[�p)ma�:��5%������;iC5PA�L@���n$<�j��Y����ԕ�3�</�	g��:A�:1�J�������m?@?�b=��<)CP�����������#����Y��U��/��u�e�V�v�$z:�$ _K�Z���_�#��YIv+�����A6�g���v�u}��Ґ�IP��FO�ػ�#:]�r��:h��z��ޡM_�<�+7ۅ�ײ����m��:�c�<G��F�^���I���WL_�ݳ�~�O������[��}P��Ȟ����k����*7]L�'���n�{��
Al2��=��Q���K��0����J�-��̉C�k_�Q����o�C�[��Oۏ�I��?������oS����Gd�>ț���V#VDoQ�Я8ST|{҆+PJ���TL��Y�*.���`���S�����)�*�,ӡo:s�ҧ	�K��d���$�QP�����ZKpK)aU 66s�]c,���{�#o�!���Iә���M�ݯ����o�7�<��k�v�ʝ�����'�w���O�m@��S����}��r/�S~���^؀�ֵ��-�C�h)�f�m����y�T_uCF�����[�~?�֗�~���(�?����>��V� @�����nz]3���_�����^��=w��9}�8�Np�͙�����!���޹��O�4,�/�d^f��z����@��O\3 ��+�!���6,�)	n��^gM�N�Y�= F�?��r�Ҩu��nnn� <*i`��h����[G̞�AYiӞ����R�dq����a���<��E�<�� �]TnzDMģ���/��>E�SՉ&�ߘuF�Q�iJ�J}UP.�z�z������Y�ɴ(�沠z��&���+iU���ՙ�<Z���S/���QW[�����tm���I6���<�Z���ܧ�Cu�֦K�����֚,��tv�&Q�G��M�rxV�����@�c~lm���D>eIY�� ��/A�9�wf���i������t���r��ʗ���S��^��X���������!��٩Z�B0�ۼ����1Ȩn�XD�	ci^ʶo�ժ������IgԜ!�?��ɂqA-���̀9�/�QO"[:�b�@���hY�9�.�̍�ZU�U��4�~omɛ�4�2�K�k�"��6���/�'n^D$M�>�2�?i~:ZP���Ｈ��D�>X��;��P}�Ǒ#{��׎g[�?�G���?�>��^�;������K���yt�Y�����C���_;��f^|�D����\����\ɜu�L�uK��g�$��+�3Q��->�|(3~�Гu>���|zU�B�G7�-�_���f������w��}�镶�y���"���2�����lI�x$=ժ����Z�0���M�����G��E� UR�N�'�m%����_�%�W�����9����#��@�q�E�ӧ(�t�L�*����R9�zԣ�GX�WiΞ=�������F{�����������!G~l��*�YVl�4;#��x��?܎�Ą|���K�}�<��e.��Xۛ��˄+k�&�2x�����	�2I���� � �Fe:��8C{�~��[���j.]kWo��<h�QN`y��4\���#��HB�o�[����󽗗��i?��g�:�ّ��h���޾j�?��²�����+eR�1�W���+A��G��n��1���G#{�Y�����_����;�i��V;|� y�n��������i?����?L~m�N��(G;�\��3+����k��e'�����$��Qc��c_W��t�r��FP4��]Fr��`�Z�e!�[��{��S�l�F K�qm��' �u�%=~nr�
�� 4٢��9�G����ʐ��(���l��<t<��rf�Fܟv�ν(*�D{�7�w��[�_}���v�О�ǵ�w�_��G�O��o����?�,���gr����P���q�L�<PH2�6�ިl䳲QW2�{���0�{�9�F�챱�����7ڷ��A��.Q/?��j����p����Ϯ��\jZ
���ڂ�X9�!؀e�/��x�e9x�`:$ߒ�AB�z�V��)����g<]��\�Z��� �HW�5)/?e b-�����U ��LP�eo:��kI�S @�*�Y� f���f��V ����K)���2�e�(G��|S�w����Ll�(�� /��d>�ү�c�:����Z���1^V�I'CYG��@��/d��8��|�����[�P�_ןykLϟ���߽���_����1��Y`B��,AhhM<�I�˴5�	��,�3� J{|=�<�F��t���O��0�9���N�2�#t����t��/eÙ���q���Nښ5�U(�F苢�vAz�+�_YYX��܆�4ƦD�5��\�c��q��/�,��9���`73Z�%�%yW��J�8�ܤ1WLx,���2��:�v�::���`�h(��[���i�l��nf�'� +>���'*����̔SF�#r=nI>���H���ʴ��$lW �8�Z�f�
]t �țM�g����cG��7^?پ��w��U{n?Ծ��?o��;��.n�����ε�}���[o�kǏ �����|�?��ڗ�=��E ��,٫6 w�D����-=���_T	<��+ ���X@�'_\�D�������v��1�����~�����}��U�;�ہc�5�'E.����Sfr���B��l6�Z*'U�!2���d�ʝeZb�V�j/�BF�t¤MF���٭+�gAr�{�:52�z���W���`Qיteu���(����J�p��;�����;����{_=����s��:XR�Z�#��Dg{"�A���pk��v���rr�맶�CR�P�)������O*?es�J��Z7�ߴ1�Q�0톺��_|Iԓ��W�ߺ����nԇM�ky���� \�GdT��=�we	:�o��/�ܸp{�=aT��՜ˀH�˔�Rf�J��Y��0����6y�dyz�������Z��U]-ff�wfvwf � i���o�����b���7|��F3�H��+ ������.]�Zg��:#3�<�soDV��˛�q��
Ǐ�����)]���P�PM����9G�DHIH�$R��C�v��܆�m�Nk��'?j7޺�\������Ͼm���W��/�ΐ��8��z�B����eٔ�h8J��_y}�Ƹ�<*�RU�M ��� ��e2�>'�pH,/2�&��&�7z�
3C��W@�{�2�#(���Z���7����J[&_.�{�����4��/�; r�~{Eء���n����8B�oM��u'�8k����umLW�\j��?i}�N�x�$e�p{3��߶���o�_���"��K��؉S��aʁƈ0stw
�%OY�s������DP%���}~�ׄX���,6-O	nǆ���]���?	n?!���_�
p��:��~A0�Pp����N=Ӫ��'�u!�(:a��26�G`Zߴ��WZ;�(`
���t���Z�S�j�&�O;/�\�,�;�=�]?qN��H>�`�<�����*�-����<���T@��g�C���T��@ �B,
!�גa;Q��Z�kW`��
�[e��5� ��|�/;մ�M��'q�E܄qSZ� R�c��x�#m,���.�������w��}W����D�5@D�:�=��i�uf����|�G���=ZJ{pk�o|/#���T���M��}P�hS�&;�/��C��-*(�viG�G� ��O���<«%����`���S]�>����u����r^���I{z�o�!��vG����	�	�����tO�~����=�A�㔲�K�G��RTmɯ-[���q��w䛪���
ܖ��K�P�7��ۼ
 �?�_���O��/���	]���pI0M�eq6�A�.��б>��`�z�L|n�c�}�`�}�I�[-�����ӧ���W�;R�Ż�'�s�mn�\!����4�u�#��v�:KɋN��i�l���M۴`]˹@��KNVv8�q�}�w��g�9���v��Ӧ۔�˭���!��f8Ll�>�sc�1�W�k� ��/Z�a��>1f5俆��}>��_A���5�K��R飌�AC���ϵ���H���������/�EV�?�����UF���Zo�C�ϑ��v��)���������W/�cG���v��6M���!U!w��29���/�%�v����k���=p�C�/�|��������s�u���E�ѿ�##����+rOá���YgP���5W�Y]��Ժ���4��wqe���7[���S
����܂���jG��������^���^ Zb�UÄ�!��7#��
�Z䰯�"�_��D!D�Q
,:lm��) )��a�������Z{��p{����j��/����c|~��/n��?����/
ܮ,/G�;60�'N@����0�óh�Zm�?Y�}��eL�����ƭ�|0�v��d|�%�V%ZX�����
�[��_�E������ԑ?�_�Ԫ�0�H���V��2)�m����R�l}���Qi��y6	]^ÈfIFҲ��%ٓ�����Ė�w�_��7�ٳ	�'������}�{��7΢8g�V�~�ɗ�׿����W�P��h��s�.���������;�8�j�Ơ�j�ZKhW�ef���Џ���:G@.zp�����?n�������o�_���ڭ[�}T �Qo��J�`'��$��S�U��D�)�z�!u�pt� �s��ݾ~η�E;�pK�lj��.���M@���b��,���A]�c���Y�7<��_�7���
��o��Zkb=�-��Ǝ��,�Oy�t�1g���Z߼Xn-_�+a%G_.���7?�Ͷ+(� ��#�}?�O}ڞ��/c��UG���@����8�������\���̽���(�U�F,q�LS�)+H����Q�x�N��?J��ۗ/����e'�ǝܮ�<���Ё!�$�~���(k�H(ꂬ>! �9�#���'��I�D��w�j�4��B�����6�(��b�~M}w���%�Y�0���i��*��QY�|W$���gu7�ݍ���=���)K��e���$!nTb&�Ϳ�{�bJ����q�S�*��Y������{�3��u���;v�YZ9��M�M"1i�b�,��&qb�h�z�l�����6<4��_h�}z����/�ܜ�r@�g 8���f�:YG�����tst+�Q0�#���K�Gn޸�h(��G^SF�͸�n	�ϝj#���sKx�l�}����O�ɿl�n?@=�د� ������<(@�m���#<���o���Kd9�7�_3ݵ��S�p�>�8�Uw��Ex��o۞�Ҹ"C�|`;�0�y��� W�*:KˎWh����U��#Zn;p�c�������g��W�٦&&�G�4&����f�FKiǣ��������
P�!=��m��#���U�:�N+y���UO�����E�i_yUZH#Jo�I��ߺ�%џ�|���F��p�f�xf\�B�JG�2�(\9(�u)Y����?����ۊ�D�i�1�s/k��V��b�A4��'�Z�f�X�PG�<��=�G��`!��32��R@lQnx�:n�pw?u-m2���x���h���H(�bs�WVp��ǻI,��~��U���w�Y������Cv�����o��[��V۸&r�Cj�F��~?\u� �q����n$�����4P{��k�U��\�Pr���6��!��$�A�2h^�s֮�����]���舓F(�`��U{�����\����e�X�N���.U�6�3������p�}����ƍk�¹ә��f��h?*� �3���:��w��u�s���dN�| _�-\F(�ܞ?M���s7=3P�"���r�NXQ�;�J���B�i�K���%�J�U'VB�ڛ��f�_��B����x�@
4��J��l�='����cU�ι6��=�J�������ݕ)� ]�ח���n	5ib�(:p�o�<$M�ѷO�+;Sˢ`pǬ�lp�z�˪�-����&���܋�Y0My�!��;�!����'�u�ݺ��5���6���SwF)T��ͫ�o=��|�~����{������/E�����2S�{�@�+<���b��RW��7�R}w���,���:I��~�;�4��w*_�	���=O��������
���ܥC�����y)�4u'M;��e�<�u�����ء�N��=ߑgS��Ĳ�#*��[`��e���TV�z�wC�$/^�_�0�u����Ϯr6���ʫr��V��%5�Z�"�����^G/�):��+���U^��o�߼�F�g� Ml��4�#s���OяF�m�驹,�����tʭ�Es������E]��W2
U��+�e�nhM؝]�=A������E��IT�4��=���JǒA��ǎ�f���W��(�����9����;�edfOg\P��W��E��m��3�mG��y��jF���NV8A��^����
`=�g*�������~�Z��������ṊC�D�öV��95��u<�{���zO��ߺ�̅s���via�=|��qV���fL��W��hr����6�6�F�]��|dW\5�y��z����G/Kr&��Ʉ�K�Owݷ�	��O>,��qU��ݪv�|#�'��Е�9W}l;�}������n �z��R�bSA��D��02lH@����hC�2`��@;���2c�@�̎��*p�0� �|-,|e�?�G�[p?�s9�Sh|�܏P%@u�u���'ڭ[����l��$� m��1�?���F#$���e"}k��j�����]r�f�K gH;)-�g2+M��V����$�n�����9ņ�
�m�&�b�V�Ͻl�'�V*v?/��S���:���3x��K�֋a���Ô���rk>�rax�mzr*�q��˗.d�#�@�v?��$2g%+ O�>ݾ�����~�KR���M��Mg9���Κa���BZb����9�i��_x��&��>9.�G���&��=G��e�,�ekf�V�Tgy�4�J���3��ֲB)>�Z��=�S�8���i'�xN0N��4j��v;C�U�4���u�>�5J��	���0�m��s	(��^3]��Z�%~��}�]��s�|;b�u-E�Y��{]%`�ޡl}�jK&�����*�v�}P���ׁBGtj	64j�8��s��� H�n;�s�=�C��	e��w=�
�/��9���u��ݍ�7������x���wË>��ql�p6tߙw�|�.=�1J��)HӁx������3�Q�:�ޏ�5�'o'�w�Ĺ� �E�p��o�)�ݪ��d^l'�2m'`�v��)%��H���2A@&�q�]�j~���Z���tͿy�wȟ��49�֪�J�I=9�'hH���9�Ew�*sx���r�_ $@�O_>ۡ���5��N3���W���R���Az:R�{�w7ז��:<��N���L(^��!�$י��%ߓo��p{0nS��x��HW�g>͇i�V���5��x0}�kn5��,���B6ZXX������i[��yM���6[}��Aks�9��s�>�-��O�a�%�?T=�+��cֺ���Y�nn�|p�`G��_nۭ��쌛=h�>�<s��L*=C������R���e&���9G{�q�6(�i�z�/}'J�m�6K=E2x݅�D��:�F}�[nԔ����o;���w��F,�ѷ��a��r��MK����#��\ld8�~ei�=y� ef)�;��>�>��k9=� ��ؔR�ȇ�
��4p�H�������^���=����3�ٝ+�"^Ƣ� �}B� >�$��ٙS,D'�=��ֳ4��%�:��8�e'�������Ϧ��[�������[n	�d-b��� ����AL3��ތ��^P�J-��K6.C�������������q�ltK8�[»��-�������7;��}������wn	K��u��{��+���?�0Ι�Ǜ[�U���▰���ڵi�T�
F�T:�-�����9���h&!iMɑ
�
�<l�|;�Ӄʩ�B���B���+h��9>���mi]S;Z8t���?Z}_B���e.�񵾶<;p��G�,qK@h�Q���=v2�h��e`fj����_�������n~{+�RN(�������~�z�l;::_�g(_|s��{��MN� |����O� {�)��=~:�~��͸�|�͝�ݠ��,W 7�=B�f2p��w��H�T�#g|lh�-��?��h&���������TfM���^�a'c]�VLwoԜ�w���CaYrMz"�=��`���*B\iH�3G,aD��(������e��	��w/��^���qHa�<�UѤӞ*?��AdA�؛��|��*�
]��4���3�K�G;5�-x�� c���^`�m:}~����4�[RҐ��7\v�P.�B{ͻ�A�١
��U�6�n$R����{���s���Rp��<���u���8"�����x�8�\`��x�rq���
�s���-c�~h�kҊ �����H���ɍ*�Z�"KzV��2J���J�s]T'��m�'�i~S6˻SfϾ'�|�~K�*��'>�䵾/���a�s�����#������G}����eB���g>���~�G}���a�xJ���[�F&���	����q��"����o�'[�z+kx�"EF�/;�n�e��c?ON�_���扢U��u� .�N���}����6<t�=}�ؾ��N��O����Џ�#i�	��Y1r��_?�Ϲ������Yx�^��Y�[�k���tO��F:H�>����81ڮ^��>����av����l���N�/��?o�o=���C�#���"���%}*��|۷׿퀌����C:�P��:JU�*��gS3X/��-W�<�I�Ю���)˂��*�#�{�2]�tH����[Zg��L�G׹Χ�xxU~7Q<M��*�qK��[��?�a�|��`o�|������gg�#O47�qE�l8����)��T��f*�J'ie��v�Y�3��U�v����u���巍E6"/��<�&^ǈ	�K��L|'-�su�q�;}o��������d������Mr&g�L���R[Z��ݫ$�,��On���?�'_�~p��p�2+��C���a֡��0�`,x�O��cZH� �a�G�/�J�c4�4�d�:k�]��-*]���Sw|���ZN�<�Ӏ^�����?����m��}�����a��������}�ClKLa�W���J�v���e����ȟB�6-�����|�IMsDQ�ȅ�⻴Rf�t�j�jF�x6���j��`ڗh�/{p���n������A�·��vfb��-�7'��������\҇1�(��~��G��ةvD��u�������o�l����_�5�=�^����O�^����o/�j��q��|y�N{���������~?[?�^,Vۢ�M̷/��p���_S�s]�Z4�Pўl�=l6�_�$/��ٻ҉�-�t��$���p�QRw��,��|�-«ΠV������R�Tr*_�����Ⱥ~5ܖ��5�N�c^�e?g��	�8m��" X!ĿԼU�;�g]���<��y�ϡ }�w��^;�+��1�.�u�H|<������~˳��l�JM�R���K�/�u�`nM�TҸ�?�����FƳq�r�;uNY |i���<q-͍3�V9��5��c�N�b������y^���w	���.@�˃�tq�`ܯ�[�v�o�n�Jmtt��K��ԛ$]������� ��L-i��c�� ��yA6�'�p��[ioκ�\�X�<�O�op�������
ҷhc�ߑf]O$?���:��u΄�JΧ9{������<[uOHr���̥�{˕ߚ�����_�&��ߋ����=��K��dI�i���?}̋m7[v�P�1��桻ʞU�5_ >K��Z���6�"m�7�T�s��� ieJ���н(QO�9vl��}�J����������gO�ڷ��m��ů����n���%�j�!&�I��x1%�2�ߺ�>�H�l�I����3�b����E }��q4�1���{���H;֦g��g�����ݹ�s9�����xL�\�7j%��Q�w�H]���r@��g�Q~	Z��D?<�U��<-f���~�\����	\BOeE�qG1�-��[��-�_*�՞d�\��Kn}��6[[_������!�PX&1Pdi�#?��p��i���L(�r�l��ĳ��K��gO����aG�P� ��F�a��O1(�ɏ��@��|��4�v�t�1�B�7�����;�G��jK�g�7:�͓�E�	]C�����k��	�VV�ꚆGۉ��Z���j������>~6ȝ��@8��ُgS��Cm��Ͼz=1�p���[���!�˥=����9�.\<�9Ӯ�� Wp�/�B��f�b����pp�w r�o������4]�U?���z�b��o����	��:�vdt�����W�*���
ܾ}�R��?�8�֭K5���Ԅ�_̤���]�p�;�� �6��gOgaqw)�E�)�d{;K}\X^�B�K�
sX�t�\{���R��ԃ�}����F��Һ�YW}���i�T��8�-�Q�a���������[��㦧?���H;z|��bi4.&?3��>�������nn�4/]������A��y��ɬI�:r��/�P���GHo�ǿ�.]<�ِuaq'�;���[wR��\�4^�5�X�w�^t�ju��:�m%޵n�Znp{^oe)�w�r���������i,[���X�&3|e\� F)«�up�:#�L~w:�i@
�,��_2�����TgPB��8�{���8�P��]�L2��ks�7�`[���|���[��{�6_�(�;^��1��^\~�C	�J+�RC�����"�����fM�|�=���s�p�J���k�#;�=��4�Y��.�=��a��{�k[�t�x�un�r�/�v�o������:���)�q�ỾPi$��|�9iu�$Tg�?��^�	��y���F�u�L"���GeS�|����7�p�����[���L]J]B�e;N#&͝#�]�����H��fVS������p�!/e�,���|�th�M+�=K[�`�ç���ş���z�׭�|9�}�Ý�|/-�#�����Q��7��y���/G�M�n��$ե�|X`��p>���9���4����sy��4J_�!\��zW�d��sH��-�7|y��">�޿t�lF��~�js4w�{��i���o۳�ɶN~7@M�N�X�][O�[.w,���䯘)1���Z������W�|���ǉ�U5ݦ IwUԝ�M�}�j;rd�>p����_���jw;p�U��aW١�L�hۭ����0]��_W��Q��*���~��+�;�9g�$�r>����z��	���m�Q��Mi��d��*�'����o�:���S�ۋOM-����� ��Y_�:Ϸ�[]��^��u)�}�.t��צ&�����m	�r��)p�H����9Y�rY_E�⥊�������YrL��|{Q������g��G�v��>�;��@����e"~��\��@�2|7<Y$����e�4 ���<������J{:1ݞ>�ȝ䯩��N���>::���_��o_O�.|�'�'�k�i18��j2��N�	d�ڋ6v|�=�^j~x#��
@O(@�D�Pu����
p��<�h�~�u�曻���'YlZ$�o�^�QhϏ���h?��ڵ�W���1 ٿj_|Y����ߴ�g���G��n�˗���G�'r�aE�J�qi�j�
��5���V ����ӑ{p<2�֡j�=!���%�z�-4���dX�J��v��*!�S�xM��z/L��E��"�vus�J�8�u�-�}��.o��h-��jc��۠G�*]�ouY`��<�h���Gi0G",��3+�&��_����0;;�N�9���O�~��>h����گ�;�dr�}��-���|b�m���N�8a"'���V���)�r���Gh_�n��	�`�K����~w��a�ة�Y�q���s��Y��X l�G�|"��|�a�ԧ�~8|k���΢���Gw6_~�%7��/*Һ�9��9�Ѧ\�z�Y��b�<��BNխ�Jv-����]���A������_R8y�s��.���;?M\�ٍ���/�Ǜ�,�r�0.S��(a�-~^��y�ƟS%`;�2��N��3��?5����ʟ�5�'�<7��E]iq������O�i��ݗr����O�pK'��}�N��5.੉"�̱\�s��Ȼ�H��"!�`\�X�ϭ��q��s��g\�K��P���q$��]��V��؉��`U���Al�"�H�L���N;��r��~ﵬVAyX�tZ�T��3?��Ǝ-���u�w�	��r�?*��[?st�v��E��)o}�Ų�.��&�F�#Qh��ݧ����C颶m���q��ڧ�ׯg��V�m�n\��|�#�	��ه�86�N��6'%o�7/.�fR����om(⤨F��O�a�K����C���[�	�Ѻ�V����$ۯ�}����"W��?e+�!r8y&Q}���ۙӧ����1R9��|r�>�^�'�ߟ�:��S���[y�v��t͑G]�(�p�X��߀������N��>x�]�X[V ��ik��пoK֭h
�C�fU���)7��)�ׂ�M��k��������S��������g�ɓɶ��S�El�[�%��׏Wp{��x�Z���ދ���}mnf�}��o���<x`4�d�e���ܺ�E�����M�'��iǹ_���^Fe{Z��|�������N�[��H�!��*�P�!�����L�+�r+��i�����e8�P����tw#p �]�ܚ���t���@w2�p�P���}
�^����_On����=y4� (.�K%�=-�0�>����������*�r6��b+׭
c�P���L<r��d�5�;�~������l�~}/[W�|�[�����KO���'�׮^���@-�K+/���r�p{�ݸv����>ȶ�����h��SG5t�m駹���5���7j��P�R����˧�6����C#��Bz�弾����u�ۗUl@���#ހ[��xic���p��{>І Ӛ�Ik�J�Xu��m��5wd�h;|���s"�
ڛ�t��  Ƈ��E��Կy	m���'��|ھ���v�޽6���r��~خ\��v����g�'���7�g2����gł�%���T{��Qv��D�R�z�M>_���G��S2�4��඄F�N��eX485p�`F�G8^�|.Y�[���������<�)��:�b��f�,��7�O�y�,���6��'��<)Gw�{E����B�o�	*%m����}V}��q�u��_��G��:�|z��Mj;��)�+�����#������g�[%ק��X<���������?;�g��C����/��+8�h�������c'ޒ�|�3Û}��~�o߉�v'N��w᱀۲p�7�ɫ��a�/�+�^ɣ�?��.��A۬�W�v�����Z�]�$�Ty<W�mۂ���Xd�c�u[�#�s�	p]���a:I�����O��A�8�b]��.n��{�x{�m"2��{��w9w�|��8�2����&V������ݹ��;����Ir�J���$q�ǳVwi^%�B��αNB�ۆn�q�7"�jߗ!띣` ri�'��Mt�飵��v�̉�f�>��H�j߅u8���5w�2
Z���ʭ�/�Ϲ) ��V�I]�}a&�I�(�#m��`V=��xٞ<]i�}v��7�����gD���r�4�����˟��W�c���K���/��^pǑv�����޸~�n����G��s�m4ś]Z��T��y�]�TpK=s�{;������4�%^��u��'��ڧ��_�i�nݏr20<l��4lúN�A?����흷���>|��?{���ϟm������U��ce���U�_�X%�WԌ72	�����Έ��`=��w-��T����M�����,�:|V�A^��V(�����44<��o:��LG�]���G�f�Q6�[E��#���/��������gm�k5�������{==��n�~�ng� h��8 0����n�O�8�gQi��v����l{��Y�hZ^Y���\S����O���{ml�D������}�~���7���r:�zk�ޏ�%�}+�8��a�k�/��_�j!��Rp��h�O�ڕ��G�'���WH�X�|j󍪑�j�U����쭍���}��F[OV�p������n�G�TSx;Ku�J�zA�`��Ś�/@��>:�m ����e�C�֑�ch�.�8Dx���ֈ��;��@/�ֵ4;�e�t�? �u�C+Y!���,ՙ��7�Q&�h������g�'�?��]�~���J�<�i���V�������;��h������������A���R�!�=���EefT��	n-N�A�����˝Ç�Wrv�k��
3>>
�=U��Sn�� q$��,�E��Z�R?vFT�!33��H�b~*Oi��͖�����З?�QF�  ��IDATj���5kd��ፃlԙH�y5��1]����)��9���0���>���Wݭ��#'�ɗg�-�]���J��W�7&�N��c�����=W��o#�	�n���Q����7u/1vQ�^̺ $@ۿU���P��"%Tɣ/vqt7s驏�S�5�5���sw�����3�\���KRL�h7�}���_�|t�y�O37yϰ�|�ў�������vފ��/U�<ʃ��ꥄ�ɟ�_��.�W��z������ /2�<���p��'����}^<r������a$;W�9�G��.���<����JJۿ��;��w��2�εG��[1�{�_���:@�>z����w�"�П�\����È�^�s��������I��@DZw{���K���0Z�'ԋ>1���˾\}�1ͺ�9�{�m^�2g��˗=|0۾��~��O?gL���0���7��Q���;��p������m��H,��w� p{)~��^�}����%���Jb�FN��9,g�(܉<�p4�#mj'.zA�>�E?���d����=��{��&`l%���C�=ܾXk#G�k�η�ߺׄ�g��}�+z<yt���GZ;�/x���1���!}��?�Ȫ0���3 ���{��ߒ�����\��N�t��x>.�׃j����$�B�,�
�m�`�#�I�5���SS��%0������5'#.����Ϟ����w�ɩ����|p���/���ۇn��;uY*�[��u��-�u;{�X����w=�{�ޣ�������险���i��fg�T�q��w���ڕ˗�Ծ���T��O�h���W��O��^�#n� ��܎��,��[-�� �4�m6;��l���}���Y���1N |4���{o�������'@��2�x��f��e��J����֗�<.g�*���I�f$���71�8�@�����,�2\���1َ�,
n����m �ֻ2��vt�8
��FB���M< ���$-0�����֡s��<�G��n�m��k�Ay��o?o�W����� n�׮\��>}6�~��;�S�/����z�t�4����|�q��|֦�'��mpx�9ю��A�:N�Ch� ��mm�	a=�MV�z�F]K��wU�//�Q�B��%=Z��d��?� �ҧ�VG�.g�Q��B�N�*u�٣�_�  7�͚��$�$�CO�ܦA�5��8� |�Hз9�H<�S_�T#���qZ}��M=/� ��\Q��`�/�^��1_�����!�e�DO�ny��b! .�W�M����Z�,u��tb�G�J���w"�̃�V|e���|��\w߽�\K��Q��3��������_B���lu��k�T����u/i��
D��zTiu眒�4A����1�x������y5���%��/�{m�Fc��1��|���=��z�|�#����~b[��7��?��b��w��g��<���s����|\ϊG^P>y��C����Lx��s��9/r�����x'���;���o<�6�EG���N�V�������s?J�~��<���y-��P
/���_V�^x�:��$Qi*.��������:�QV�Hg�hU݃���)�x�0����������u�q�~���uw��]>OԜßy�w+B��+��ꫬ�0y8�n�zھ��N��\�mW�ჽ��`:�V����-�w�7g��h��z� x��Xp��������~���++�m���B@�� ��鑺ɥ!Z��9e]���� "�рE�a����Z��������g�������/�<X���c�T��-�hXsi�ё���B{���XoϞkC�&[���1�]�2��ٶn�.9�E�G^�l3����Y)jKwB}��#���a����x��Q]�y�m�Xa��y����G��+��T'�>:Ԏ�Gǎs�`�E��?=9�f�]��5�`<p4�#�":3������y�=~����?�b���_�	��%�}<�f&�T|��/����%�^g�޻��I\�����o�D>m�����c��F,��>q���{���w����w��P����W?����o���,�/7�ѡ���n�]��B-���l�~z������7 �U���pܞi?������u%���OY�JRu�����:g�n���e�Ou�4��&9���<
f��Hę
-��ڂ�N��8�ЧDp�!��u��������J�����F ��@GE˝� ����<��_��6np�2i:1E�aC��޾��}���
�?��о����X��*���/�O?��w?kK+�����V��|���gШ�#\l�#c��<����>{6S�V�²�RCZ��d�\�PW��bA)(�t����������� ��&v�ɝ�n�H��E\�C����oV� �gx�����<C���K{脚JS�p����=�E�N�f�Jӌ�84�|��ө;[\?�J���w�x�4�X!�����i�G�ɋ���Ry�5���X|�X�ʏ�s����{^�М��A$,����ߙs��0����nyy�c~�ӶE˷����8���L/sm<V|�I���7�WH��(v-#n�l=��?��Zw�#�ǈ*`���Dj��Y�ݐ��#�I�w����V�9 W���
|MB�|c>����#e����?��G��s��d�̟�su�[t�:]�<U�ɗ�*�J��/ݍ��}i"�[��o���^��w��Or��.y�z�N�:ϳ��$nB��Է��eH9�w���u孮����9o���j"sY	���_/�64�����E�C38d���A�`��e%5�g�hU,�����?Ʉ�N!*_6������}Y��˪����g�b�+}#�ڮ���Wm%��ĳ����\[Z��=�dRp��I�u�g���<|G�s�h��u�Wϟo����'p{�"�rOF{�<zޞ=������� �� E�B��X��?��#��ޤE����O'ĽxI��7ns||t�]8s��M;|�p��p��f�"KY	n�dix
���\�{t�H�q�B�q� �==>� �o�������XW>��l�t�����С# �!�?u���э�u����^�~J��A��:��ͣn֫4���+z�F�9���A-����ۣ�F�ة���S[[`�%��l�xk|�^�6��K��353�n߹��=x�����\���_�ۛ�����%l�0���9����W������Wc"��)η��l~N���=�ƙ�2��ԵR?����o�[�V{뭷�\��g?���[­����!���Xn#��KOǽ�,��$���
�Q����������H���[��{��5叝8F9D3ݎ�H��jx�*�7L�6��!'��������q�Q��*��>~'S�v�h���/���8���P �DZf\|{mk�-�Ѣln;�O-̸mo�brt�hhh���m"��.*�=��p��ӭ|,��MNε/���>���W���t���8���L(�������O�*�m���o���l?���6;?і����j�R'�ml�����cqK�ή�n��4(�琘���W�|��v o�O�	ٸ�
:!\H_���K:���W#� ��U�X�.�4��MoG�����|��-Zg
"iggdHg�O�v8f�+J"x�ȭ>_^�ܸ��S���෠I���Ƀ���^hD�}�J���+(tx��J+y$��5��=יHaY��=C���]��	}�M����5!y2�u$-?���7/�y�<{Nd��(zH��w~�]�5��stߤ��C��?�ny�����V����n~�x��C+H�[�ƨ�9?��*bGV����J�Х�z^K�S-�Qg��+���^�랯��)˟*`�C)t�D�/�y&�mG/�p�rpp;����;��޶�y���ƶV�+~H��"�\�PE�J�#ȯ���kn+��0.�W�H�N���F޹H^9~�y��.]z����A>|Ï*�������y��7�͛�o�i�����A��c�g�h�Ҿ!<�q�L�;�˵9�b�0�ֿyR桄J�3^�S�d9l��E��_���:�����$c�/�A�7��v��yn�<>�WR�ę%3B�5|�����Yi��Z���1x,jW�^����'�i�%�X8Lo�Ǜ�o�ܾC�6Hs1n	�'c�ٟ�]����֙����o�o�=I�{���6>>��\�hY"U7�O՝���l����܈A�M�@�S'O��~��$^�}�p���_j���}��W�C �C ��$ָ$���v ������g�ɱ��<��m�_ P�����AB�j��o����M]e��U'm�B����-�d�ޯ���t3��������N��AI�x���ϟeT(%AE2�H[׌��C��ɱ�ե=�S��0�؞k���o�������,V:��&�G���w�_��JO�=��?����\7���!��4�����^�S�#��~�÷��>z7{Y?6���{ؾ����i�B���v�VW9�r�b���}��>}�J��M�_���9 ��o�	e��rc������A��$�V�����.eF��vzf�}�٭��o�����'���Ï>.���3�, �֜��k;t)��0D�H�P67=ݞ=zжp���pb�DF��Z�D��c�h��H|2>�i�5#�A�`��ހ��.	ˋm�]eh
SQp��������k��w�p�4��6���j�j;�`�}�SFStY&��sӃ������}��ܹ�e22��eB��B8yEp���O�'����◿n�����Y4�#{a�%�|H�4�����x�G��WV��J����T؉��.��o�wξ˵��Ne�F���K
Ct��[��(U/��s[��C��7���QN|E����C�絠A�n���w>vv�vN)��p6O9w����SGw�����ߐ�Đ�;�ʿ�^9�<O�W�*X���G���>�f<��$��b��X�������K��=©>�'$�o�>  i�����Iz7���w�#GY�,o�[�W���T���LjB�i��Ǻ��~_y�'\za����;�f�أ>�[��[�g^�y�F�M\��2�?�Z��&-ޱ�٩M��_ױ�x�O"�9B��R�Q�9��JIx�Rz�)|nD��^QFvi��NrD�+A�L�x�at�Viݢ���]��}}�����
����N\9�xr��u�~�w�>�G/q�����?[vi�]���a#�0.>+�3��j����U�i�*�D �x�s�gN�3g��-�W���yѲ�Oꬂ�G�y)D��$���b�K�?e�G�t��C�M�(�	c��n��捈�<��_����pH����z
rm�w�e��d$�r����=����/�IORw�� [���9�d<����7|琪ҧvP�_umu>n	��������?�#��E^}ݞ=�h���o��_�l>�U�G?��v��E ��(���}붖ZA�� ��Gi�(]��=�D_��ɣ����¯��3g����G�υ��?o������W_�/����W�&�se
�
Ip������o_n��/]8��ǜ���>�Ue��tb����o���::r�V"=�zr�L�1�^�2rֱ�˥�Kc��RW��Փ#/�/�$}�<`[Q�Aی�ç�Q1��G�M�[�Ee�>�8܆�"C���a .
���q�MML�����,߽n#GG�e28�aq�ݺs����lO ©���_�6�%����(����ӡ�n���l'���������h$'�ge�!����Ҳ_��i��!huY�/ ���5�����g߶[�
KK�\�����<�._B�����~P�������٭����/��~�
:xp_;}r��u�\����>x�J��=vl$�	���6�0"E��4����!�D�x��^�3�O��'O���WX�6X�R#���y�ƭ{��Q�ɻ^G(v�e"E����k0�B��� j���]m���C�u˛������ۡ�0/c�V{��T��g�4r�a||I����W^d2�?���,>��������]B#�
�O.�Ͼx�~�ɷ��?���X&/(7/Pt��W��L�އE��i\��� x���pu�eG����(Z*��{9x6�[�`q��\�<�Gxe]>���4�@]d���pz��zN�F��no+)�1�qxK���z{��΂�T��<|��l�~��rĪY��4l���s��u�k~�d�r�<�
���w��_�I�>�C[ig����<��V׀��ܱ,�Q}�;�BOajǝM�c�ŵ�ų9{�jL;�� t��y"!����D����j��#����A��f��.M�J��hz:�Ho'}�������%vkLwJLޣ�Z0���W��Ȗo<��<�~�{~#��c\�Q��;����uT�*�ռ�vܫ�au��9��|e�U��N,�k�/*J'��U���ؓǞO�s��"�"Mzp�K��7�?�y�[��n�+60���s�O	�����c��TZ���j� �'o/��ûNp�w ��dǵ~�?��o^�M�x��`�DȎV1n�A��M��Rp�̯��(�'ivu��y�*�B/�yϻ]��v+,�U��>�}�`�k�ǌ��ϲK��2t��GIҼ�f�U���J>��|՗-�|T!�]}�<���K�ցC�~�'�s~m�;�2�c���	p-��`�(�͏���˻|�%�);7̍mW�Z�*ch��w� �6Z�5MG kU!��A�;t���G��#�,�{�T�˝�9���C޶��A��j���ЁX=��ڿ��خn�� �?��/ڗ�p{l�x�{��7��A�#,D_�A����ګ���ʍ^a����W�I?���s�f���&/څsg��ݟ���/P������?����W_������� ��Pn_���z{�b�~�8���t;�D��ѡC���Pv�s[��M�8�_�c�跲!y��5"�#a_����J,�뼛��E�z��������%렯�7�����B��ڇI�]p[�Z��Y���f���O9�|ح��� �Q����6�87צ'���g���F;t�P;:2
F;�W���q�?�Y�{�a&��������/.�9L��V� �t,�Xd\�4��>�=�G�2l?Df\$y|l���=s��;{��;g�p>{�y�خ�۷���7p�&�D˯@�0p��h�?�ؘ���h�ϟ�{ ��	��Ӧ���n������B�ui]���Ooǎ��i;��JB	~51;�ߠ�fg�2@s��G���In.+!H7�#Y��Ryҩ���S����n!,�h��ZouM ,n7j0�6�sq�e5��ߥ�
C:-���t���K䣝AMZ�-�nQ���[i̿��/h��p'O���ׯ���B7R6n�11���2�?~�V��2�Q �?��Y�r�49�V�ϋ�����;�èP����$j��G���J��/�>�����E���
 w�Sg�m�'Br�����kӷْҔ�����]�i 4�-!`��l��7o�5�=�:�d��5VK��n}����C.�t��n�Nx���:�^�т�7�)�m�dK�)@�N��?�<�C�O���[�
����J"!�O��8�D%�sg��;֫�١��ɇ[I�R��f<���y��k�rOvF5�n�Ew�M� �H��Ѿ��C
O����=hd�$��ٺ�W����i���Gy@}��}_+����W�������g�!�TK����b�o��Nɑw�C�-�L�ez���&��q��VG�r͟��UGUWr�,�0.�@zsC`C(ڗ�t?�۝�eǳ�a�S �����>�|���[�������<��PNR�2���9���^��K@�ݡ|O<���j�� �TGb�w��ö\[]ʛ�FQ����yx����v�8I��Fːy�q�B\�P�u��9D��s�׷��۝���;����L�HM�*x�;�&�K�׶{ް��9e$�:��[�U8r6o���s��۔7�g^et���	�Nv4�?���o���6�°E_d�i�UVd"�V���R[G�o"WSfwL_K��_\�z�h�&tx\�ϑu^GP�4���v�#>O��6]np�e���}��в��b��w�x�u�w�\�}�rR�qv�[��Q?~����8*�ӎ����+i+��~Ҧ�����M�L���w��J���k?�	��?<,�4"�ʖ�݉qpɹS�nv`V�~p�A{�|�-��0�����ud�@�l�'on�BK]3�]�a�+��+W�����s�YT��mq/_���n�������ms?qD.�/��z����t-�/�Fd�y�O��v�)�}��Fսёl���p']��<�V�`ve��;Zy�'�-YZ�ȌJ�(�TP�����:��������G�[7�%����<z�&��Q�H���n"�����g)=����0H��
]� )�Vw��b��W��g�Q(����{����̴gϞ��������p�FӨd������uY+���Z{�d�ݻ��ݿ��M<��[;*!ʇ��YbK\:�X�lxot
�SB��"�٫ƭVk|dmL˓
@��@�+`_tBaB��� njG��Ch<���D��l���m��u�F�`�	v���[��������K_Ұ_��m������zmfߢ��#� ��K6ȯ�r�弑-�V�k��5��I"����
Z�X�t��;���i�xb�F����_JGyA�C�4@�"�]cQ%Cm)��p��>�+,�<�ۦ���
�G��eL8b��d#g� %�# 3�&<�R5��s�>H8��G��?d�
��{kA��Z��'��!�Σ3>�V.�rW�W >���G�opb�@n?ׂ�l���,�@�x�P4�A�l���<�����V��@� Q�S�i:ב6��" `�[a �Ԋ_��t�5��k�e=B�
>ש��摼�O�@V%��*�O���g�۹�'�[����S������v��X����{��p;5~,+��)"���zw��m��@�916L]��xM�N����v
E�J�Y�J�GGG���O0�)�E�����GG����q�̹�-.����s�SH\�O���k�r�k��}���8��
x
%P�Y� �A��m�W�Li!���9g�	 8��<pX��,�ՆxE�|��v'�3Nw����NAE�� ��Ю-�X�5�L[H����7|�	��B�4���H�ʏa��]��'��֦r��JY�#��lyK�X�PI�:�6)/��҇?Q�L�v�}�u[Z]o^�;�e���6�"����Yw���p�N/�"ʾ�W�-�+;�(�ͶF�,�=�_#�m�:y�����(�"�n�uGI2�N�/��/��>�mN�h;dR&�Af<�¹����Άw�t��>�0�<X�V��Qd5u_ ^�P�1#�?Ҏ2���k&�Z^�	&�m�2�Yg}GY�2��1���ܫe�N�By�g�E�9�����9z0�ʧ�\�H�2r��x�w����J����5��PfCյy1'�M�9q�
�
�&A?������p풖�K�[����,�*֙<�
K~�$5�ܷ�h�x�]�P����'��;`���#O0.��&��uFy��
��_7�BMH^p%#���m��b����]��P�0���U]�&���u�W��빛xKn��<�}F6�g��:�P�6� z ��z��QT�^w@�d���� �F�!S��}�֟��Q޵O;6B_�o28����7����]i�h.�k�]�!~d@��"���Ş=v& C���������Q۵�fg���2�����F��[FK�inx����T��q���B�p���}�tѸ�HO��ϴ��g�ݺ���=���� `c�v����>y�߀S�LO�5A^r��ʯ���䀸�WQ�wǐ�ё6r\?R'�9�)x�b;%�!7-�Z.���w)O5q��}�+�]r� �n/���\��Τ���ft=ۃ���HÝɴ����<(�*�̷�9ĢlgBe���ƫ�4��o�<Z��<6v�]�q��9s�0�������4��S>x˱|`�gI7gX�!n��Zi�W�K���Ck�D��'�SN�qZ'�P�C�2���8u<<<H����k��a?-���f]zN z���c���ԵZ�'�h�RF��WN6К��:�H���m��t�MZ�K�"��5A�[6�j`�!�;:�[.t���<\;ږ#�V
�v4����4ס�B \C0�0 3�\�]��oC���N�@M�O�����#@К+�c����^:=��_�=��6񙮀��ȑ6�Μ�^tT�$�lZ\��N��e7�#�����v��̙��(�ZV�������^�C��&!�����۶~���v��v��yd����&�(��U)�X!�r�@u�Me�ѣ.��2@>���:���T�6��*�4�wm_)�Y6��~T(��.)Nb���
�����ZK��|$ք�񉝨�h���F���e��~��Z��/���@]��?A��։nAt�k���
9q�)d5�O�-(��q��z��U�x��(��%�&�-%Z,�Cu��|G��o╩�e�3�Ë��a��"��В�x���Kd,� ����Eɂv*cQ�ho�6w|@Fy̖i�
�i��IGik;
��-h�jhY���FM�h�w�K[�.ɣrÑ���\q�u�'7?�@��S�����АL٩?�[��&�G��	3d�1=74����s/h�k���ud�x�u�ģ�%� ��9ʶ2 ("yU�&�|Wu=,���3�N9���_�n�����7��S����{�Ey#��,�������H�<��F��L,Ӌ�.���k�#��������%���o;?α������iCqVn]�t�~c��[���<�_�h33s�ݺQ���
F������>QBl�5C��2�l��sjr*��ϟ=m++ˡ���c����<����R�<y2�&'g2���gF�B��#K�N��8ʿk�*Kݨ*�G�R��M����Zˬ�Ĥ��V_bw/S&��*7�k�@�6l0j�9�����Ϫ�R�����y�����|�[����ri����72���U\�Rw
ۥ�PFZ�ꈆ|648�>Y�T�baa1[���������[@���j�ZX_����wB&�a���.��6"5������LNMgS�9�g��Vʛ���^XXΖ�O�M�Ph9�hf:�]�:(��E�-c'��Rs�z��p�6��ʋ�lb�ݾ� ��%�F=B�z���:A��Ԓm���)���6h��J�͔mXN��R|b��n_Z�_�Ϸ��+W���  Xu�Q�\W��=c���>����\k�a���Z�onv�N?8��;�'�����r&8L�o������5#]����簓�)g�WW6ip���[m~a!uzA+�u�!�-u���&�}$�]^��94Y��]�݀��/i(C?�ˀ2�$V�b^i\|o�TʑBU�Br�̉v�ܩ�K,0P�n���?���7߸����c ���^������ɀ��Էk��� r��vnq_�R�b�〩K��"�ƣ��9a�4F��N�C��E�U8��?\2F���[K�#UR�M'��)"T��`Z:�A4�}��C_�O��R!��}�:��hh��wn!i�*#q١c1	]Z;t�@ V�Q�}� ء����Ԇ��]�
��!pLieR�< �r�|�rE��3n�7����?�֖�(�9���Э���
�e��"���]�x�>;�>=Z�k�����۵���k��TҒ?t7���j�؈�VYzl��©������3�|w�z$�Z��E�+��@�c�\�٭���6�W<G�P�?#�\l��c}	�
4	` {�Ǎ�|J;#�V�
��»���ax�ĉQ�H����|Q.�B[ W�*4�.����2�U��n4c�`G�C@��~V�T���u�ײ�o�۩���S�`DF|�,j�P�q��2j�v�C�o����u)�ǆ���H;A��z �_۳VcA��ʥVȣ�����ˈa ��F�M]֩�5i@kۋu`�*O����� ����b�%�a�Ax�re�غ6H�X�y?`�x����?�'���R%x��!�ʉW�A몆�&�pn�iځ��?ۡ�����������s�,�'�+��e��Oq��Z۶���u8i�F1TƝ;y: ٍ��Q�(�zRN�׀���.�o� ����zց�2�L h����1�n��V��'��r<�̅�5$��j����=����j����QN�!(;��^)����
�K�T��:,�������-���N����jj���i�;��ҿ\�\��On>����L_�#���G�R�9��P��$�CL!@PMLL&8���A��dt�u������-��ۧO'��m`�!+ui���
�BQ�y��+GŠ#�wGEJp�Q=�-X@����g:!˾pph8Yv�X��r�ޑ��](���8��*��X������J��������o��2�t7���*��\�HcC�[:�臭o �77tqE/x���i���r��ss�����ר�ť� R�1���3�L�Q`Ze��>,��`Up�o�Qis����Y3n�� !2�"3�UP��FG4�]�"\����G��TM�C��p{�Ćh���a<�xZY�&��y���b��ڶ��B�3䱄� �4\�Zp�
(s�~U��LK�j�j�B�Wk�X�Ц^��G��<q�g��3�}eֽs�RN�-�@T�^��&���u������f[ἶ@ ��+�K@���߂A�"2�Vځ��[:�= ���P�W-�P��	t��׊�7粼����v��g4�{���0�q����S�pK��ˀ[}nO��4�����2"�L�U����^K�K�W/d��mCm;r�ᗂ :sj�Y�z:�y��v��e�'B�Ndk0������N��i7޾��~�Z���5 �h�N��sѲw
a=���TK���E��P~i�{�] ������g�1;��������* �
��%�z�o/���
&�u��ONKmj����ۮ�ֆo{���-��y��q�4R������H���v�����8�s|L�=�]�j:vtn�lGd�� tC�-�C��R`a��uJ��*mW�R!p�q�R{��n�w޹��_�	h-�-w��g�r�ٙ
r]��4�/\<��^Y]@���c�I���{7�{�ߠ.������O�o~�>��@O��.�g�6�Z�v�+ZXt� �K��Ŭr���ҧɳVd��J�D
e��:�.\��ΝI��-����2t[%_{ȇ@�T�K?�(j�i� h���;�wo���|u�ʅ�g��^˘���ǏrN�����=����7޺^�j�*��+�s�<B ���Gﴏ��~�o����g�1ҏCl�Z~�t�G�Q������w�[��K��GV��J���I���o�V��g�z ��~�2���T������@�x�L��/^<�}�}�	0��o�+ʳ��[����}��=�%���?|T7
�1���.S�%S��'�55�'�;�;E}����@ޕPT��OܘF�'ς�-g�o:	w#�ֲL>��{֝���ѽ#�!MG/\8ui&�j�M�G}P%��sȊ��������K(p7޺�>������ŏ�a��h��)�Td��e4���o���{Y�V�N[0~�#����J}�s�w�~�R�Ҙ��8�2�-GTJ��K�Vq��W��C��@BK]�|��1o����+y7��r����j���VV"ߕM�����~���������S����
�I_B;D���p��b��� ��a�B���ܯQG'�Zh�;�Yn�+�ƿ}��q|n5�ٟ	��� ��ʒ�\��(k��{�$�W��F�>7�ОM<O\n�$�иvYq�"�ԃhvv�=z��x*F@�m-j�a)ȿPD�~E��i�a��s^�*ɇ#.�R�k�,�:~�8
�1������ Fs�+��*��-Ir����G)����c�����EY���=q@0}[��.OI$��R�M=Sш���C;��Fd���|pK���{�LU�t]���������,� ��ˤc#�\F�YdZ��e���"�j"t;v�@�l����\��JͶjCC�>L|{��� ��ZK-[,%h,�ءܞ:y,�t1�
��W����\�{�!Z�\
��\�����q-q4dgE��n�E�5țEc�YX ��%��}a-���|M<� ����Z��wc�D��.������gܛ����VCX@���J�#MW0]���2 xE�,0�i��G���TH�LHئ�r�0�r`�ī��I@e����X���$ ��d���4�g��'��J���q:��NZ��%[Y�@�\����p���ci�� �����v�j�Zi+ ���mVJ���5�"ۯ��*|�]�A����K?L���X�!i!�;;0���}��G��R��̤��ڱ q����8�R�����zm��eO��� �t2���v~AZ�+0;w����v�sl��s����������om-�m\՝e,pK�Ã�O��[��Z��J+��(�9	B���ԭ÷�����vh�g��|��N\p��aY�ח|��N4�#����je���h�������"R�e������h�Qlq��E���X�;�jLǢ���i�Y\�˺�33�y'�Í�t:���C�*Z���`+C������5PW���N|�	���@�x)`$��k�tki�"�,���P(7.^��7*H�
WwZ���]wI�
�;Z�]5D�$_��?���ls��4`M_c�5!�6�����x�y�r���p�4�x��Ay�t��"����7 <�{� ҥ3 W�mf:G�A+�E˓�V�.��z�"�	��Ux��;��RV�Gz���3�.kk+m~nY�B�@���gϞ�W!���*��q���
�V>�*J�R���r�Q�~�څ*CxX�M+�. �bHq�_��"�b�kJ)5zp����#)����>�kʤL� �ԵE�v:8b`�
J���J�wAګ�h��ܫi
���G�9@刓�J��n�P� �ؘ��oyVY9�|���W֟�(�t���k]7�>p����|$�V�(*'T��N��(���{T��LUJ��gB�y�N����G����I��d���0�]�U� k��W1�`>��^U��u�%��!��Ek�����KԓJ�+�fTS!�_R��1�V!o�.|��G�[$f��{��!r�������p�-�� G�����In7x��I�x>�������{��R��c�j΃ԫmf ��õ#t��.-�\�q�@����qd ��<|(R\�%=� ���}vvEߡ$$��9o��e��\�by��R�,�~��p�K{eҗ7\��-h]CW47;K���	�B��I��� X�y�e�S�׹>�f�^��~�X��r��(��5�8G$���Q Wp[��	��਒�h�:]�$�#�N0�ά�n4���HK6��_�@^p���$���v�v%��a>�Gc�$�̒�C��Zrd�K�K��@��p��!hO���g۩3�s�s��䲈�y4@�C��pʛ���T��!��\��5ɟ�8�c�����ٞ=�i�o��j	�QH�T6��!'������6=������ԡW �Id�Ď�F���n����B{�|�=~2�۞>��0�s���r~J�O�O�'h`x61Ӧ �� a�)fH��1x�P���||��`tA��gf�a��>����\u��ն���8���8&�lLZ�סa&�Qg�Z��V%e^0M�S���3�B��q���@���ke��n���z�a��Ǻ��Kq40�֨@�Z�@-�-p��
}�R� �vZZ��#�p�l�k�~�j@�V-��tnv�	�9�.���. 8?�ཛྷ��R��TH�U���(�	�y�r?�����'|sÕ��[;��c%h�����~�
�sC-����7[w�e�ռ��j�Q�/�_��\e�-����\4Κ���!Q�e��+�� @� ���ʛ3�]c�5@�㐪����>|�r�������P:{֡��//�h�H�Z��t�ך�����g ����]`���,�=������,�~�a��Ǐ���&l��f��ĳ� �%d���԰���� ڣV&��t��sm>�i)T�p8�ND9 �5.((�:�'��"�mZ3Z�.k��i�/�Yv�Z�&�IU� .�ˤ��
�6m�B�ܹs����໦�`Hו�:\M����fyg��B������ Z�R���aQ^�(�Y�[�������n/��!���P�7�H]�Z���R�}Q���� ��E��.��Ց�sױtA���j�V�pd��Q��Q�a��8�h�8h�}������i/������"/FT��}��ٴ���Eڝ�}/����9=�
���Eop��k(�7 {��r��XB,� ,�W��k5��X~��{�"�[�
�
^��-�Ay.�t��wߎ��oU�fg���9�|]�~%V�P�`�	=>|��*�[]7T����e�z��Q�Z��EOe\���{Wc�q�m�c����[�C�'w�GG�NUN�GٕB�*��i�}�.urŗ�Iw�݄������������9/�ϷUڶmT�z�2r�m�\h��K;>y� |��V��?~:]�͡��׎�h	s��"���;*t������L҄oͷmV�mee)�"oS^݉�Z�G�mwN�ե�88�A?W$p�2 ���k�K����ÿ)�-��D5���hP9��`�}�<~ڹ̦�����H�f�;�@�i�f�(�\y@_Ve�F��ˡ
����'T������.��ϑ��po��~ݽ?�F�:�U�[K?�2�*8�=����!V[y��ä_W>:oJ`�T�@Bâ��N>�����*�˂�Y����o�_���������Y�6 ��{0�����wV
i�Y��ϕ9��n�퉵�wa�]��Γ�ܪٯ�i)O�o�;����'~�r����/�}�����2 FwqE��
���Rx5��t�,�'ƎQqT���6`d�����ct�:*�-��b��+����Q�*3�C�Zo�m:�pT�t9��j�]Yy�����>D����W�PӼe��:11 ��)@MM�`�/��e#s#�X�*� C�N~sS�� �I���w��2dS^�s��st���i,ſxj�@��{������<] ��V`;�}5J��"�xw~j�-Lh���fyWpk��b�B������tA��<k�[�3C�s\� D�?F9�~��ɀ[�����K�n�δG���r+(��b|�R����U�r��Ƚ0*2֭� �S��]�v�]����t�J �x#-�Q��i�458�����>�
F���z����mG���>�K���i� �z��ƚ���*ر�ˇ*���(���2�oE�P����L������J[��rq�[��^�j��	����^8�=:�%d\/�I�A݂U��^\���%�/���Z:;}
�l�:R��@@��I�>��Z7�:@A����0�-�B�&���ͯo�Y@;p�����}k�����vw��ޝ��f:�A�R@j砬�
���"����h��Q�E@��������q�V�k��	�����a�=y��ڳ6�u(�r	���ti(� ��/�aK��?�0�%Y�k6ua��	Z�r@"�����1:Wz�:\�C!��Y�xpi�Ϫ��SS; W -Xs؅��������-�|���q ��y�!i'�������G&���:���λ(!���g�9ݪ�ӎ|�w�mH�3J.������߱<]ɜ+!/:*P��!OH�|��������ĵD��e��Π�N�uߑ�{�����~��zQ2CN��+륻
����g�!��sU~�C-
���أU�}ȥ�Z�)?@A���h)߼�T 1�#���XZ�f>~�9<I}��׵��J]=G_U;Y���n}{'rS�����Q��c� ڞ���u��`�����Z����>���ї�� �?˒>��M��پb�J|Z�}�b8L�8�.9g�YF�k�P.�ĻR��gsG��!]���h_�;�F�m]$o���@���ɉv��]�[�,�*����'�3e�ufp\��ɞ��g}:��׮��Qy�����# �S�*����mԍm�~eD�sm�o�6b0����|�XqA���.�M��٣ R]q�+�]�U�Z� ȷ���ug2?Zn��F��Q�~|�)O���Ӹ%�[�-�Y)���T'ᯮm�Ǽ�;td }��IGNg�y�x���r+��_�}רW��������C#�Q۝�P��I�CyV+L���h��A�T�ة��<:wK����	e=)���:`+]��~)C�+T����/X�Z`�⩐���U�z�m�ve��ݳ��Y��#���9J�zI[�o��s�!�:ʎ�������}�����K %��E�6�|D�3��:��Ђ`D��|v&6�,��y���и�J�-a]�[�
q�=.mD�ь��^�Q�)57�8� ;F#�q]P(;�L��\�A�"�l~}]��,�Ɨ� ��b�Zv�oy�l"�V<CS{>�P��pԼb�ɵ5�����o�۷�G7ͽY��@i~N!S vqiA���<�����Y�f�R��Ԫ��94`�� <p���y�E�M��St���g� w��0Ȟ!/�����<��؀X�����
$UX�R�[������q�ߍ1A`;4�<ϟ/�-!��-�N��\|/{
����#�j�Zp���[�!�u�,�D�Aa�BP��N_S��L"2�^�ۭ�V��}��֯
�W_�lw�:�������h����Jv�����Tǵ�����w0�y���Q�3t,�
#Ҹ{�a��!i=Iݿ~}�;�P�n�T𮊖��AyQj���0�
ܫ͓ �3���q���^E�ji7�vZ�5��^�N��Q��^��k1J���*� *��K:8�w��^�ô=�}��K�4���S:�z.�ܢ�������t�
N�c?��{�ө!�_~�u���o����E�Sk�u��@�ʲ�g�2i��Qި7�
~A�������|��v�$F���ݎ���Gq���Ĭ���^���Ņ�=��ǶC�	j���;�5�xG���^9�5�e:&�^˾��kԣ����Ξ��q���M����� r�_A�C�G	�H�}ۑ�DP�q��	�;B~���Ó�{s�v����>�Z��V�S�'���78�Y�\� ߺL�mm�/Hs~�W޼ie�&��n�L=����Vv�L��5��Ve����{�k9��z��[�G�PW�ٗ�u~ H걠�gZ��ǫN�EIv�t�k������0�����R{p�i��� ����	�vX�Νo�P�.§ W����Ϩ�<mOYSF�#(���YOZ��`�Vi�w��D��4�Cp������������1$�V%��8��$�Q�
��e���e�n=�6���wo�
��U.j�{��}���٧_B�I��J�3��t������P4E�J����{�n�z�n��g1���^��eYO?�D���@��ֳViGm�a��`vv�t���[�ն�ۂ��Z6]^Peyö��  U�>;��n޾/?/�C�qR�}�u�J{Pٱ,�w-�1���Snjp�ݽ�(k�/,��OaˀZ����S9�,8@��ʊ�A{J���دx�>��'��;*�S��e�U�λ��>���Y?YG���~$r_-��g>p�N��K]�^�A�Vۜ��m�~���Ֆ4�i@ҥM��<���#0��;�*�3�dg���p���!�.�Bt�He�Q����o��>PP��Y呓��Y]�N�:�tX:�L�~�~%v�P�*�\�!���V �ЃW�>���܃�ݳ����Q�������#�<[$mc�Yːy��G^w�ք���#�u�5��7�g�w~��8����̔�F��f�D�0P�P������D�:�J��������@C�i�[�q������T枤C�2�cH��/�ٴ��Ud�s���r�}� 7� os�w$��Jt����Oі����H0jO��L�{�s {��s:@��I� �"p�'�Z[�����e@�䕕m���!h�B�!l�]d�l�|b��kv�	�FP=<՞��'�䣩6Axf�?k��>Nx|�I{Lޞ&_<'oϞLŪ��1<�|�ŭ�(ZK&���e�C��2L�T�������G�+�޴B�����(���<�s?�K��9�����j9Ѫhǫ�lüX�u���X�LZ�l�g
[��X��ɹ���]~Nlw}�쳻t��L&]�A����W�g	�T�y���qܹ��݇T��
/�U��vj��V2/߽�pw�ݾ��:��@�nj��tQ�Y:٨KH(<�s�*<�ྜྷ�t�~y�	+	�V��ꐳ~�1�$�ĉ�?�ݏ���~�Q�&�Р��~������ps����޻��˧�88�� _�޴'ˬ�Q�r�I�����G� Mq^`�F�?�`ٳ�"4���#�v2�9:ݷ��8�Z+���
��\�@5�� ����ٶU����(D B1�X<YV�e�ZU�YȨF)0S���x��L
S�z-�ߥv��c|���흷�Ƃ5��t�ɟo#�������2[�ըE�	&��:�q; e��*ѿ����?�$�����Q?�}������_�@M�D !h��	��?�>���,s�5mV�yʬ���F��0�mne@7�qV�3=�Z�T�3�_鷻��N�"�z ���9�����}�Nfu��*/Lˇ�����;j2}�y�2�k�� ��*3*���_���=��$�c��Q�`١Q�}C;���/ۗ(b�l;:e�C��Wj|х���p���-R���'˝�<��t�*D(�0��Qwn݇ΏᝅX��qո\#.]$N��j�\@�?�߻��|�}�����'ߒo��;��εp�3G#N�N�>���a��}������y�.N��5h���:���2��*F��su�r�c7孓�ƝD�����.�\vŅ�ͺ�8�ꨀnn��������_����IQ��-����,�.
�׌��k*Y9�����C��92D��+(��E�ڧ;��O%E*���������"x��%��#\@�m'���Fpd�=T
u�q�)K�!s5
�6U�U��@�{�#�:8"54t���#ۜ$fr��R%ԥBI���7���w��K�4ۯ#��]��I��g�|e"2�MS����g���=���O��y�-�r��:�~o�����2"�o�C�O>�>T|	����kԾ���.N�هD������Р���?/���vú�8Ҷ?����I�G�t�/�S��&2��'���h����Ͼ��~��/�_�����_~�~��oۯ~U�׿����7_%|���4P�Q��5�B�V��-h�l�c�v��gB�;5��ZJe����!�ܵˡfw���2�2e����Ӣ{�T�ߗ_�0�= gq^�GW�2aHM I*�ҁ�Nj��ڃ0r;Hy�[:������Ƿ��Z�:���~�sKmi��ya����B� �'覰��V~�<SS���s�$8�އ�w�H��ãY����iY�b�*0]i?t tX2|?Tf���'��s_=��:gy��}�a�Q���b`��
��H{fv�:�������l_}�%`�I:,��\��F.���Z�QP�<=�	�Hu=b����	��8��?k_|�J�S���d�zw��I4�[w�O�?��o���ۧ�~ݾ��V:�������G�Ϟv������1A�r���׿n��?���=}�$�v�uMYM�&T��Z�j�&Nz��{e2�ٹgc��\�" y��0��~�S�����}@������6��:��-�A�k:�} �C���������{＝��sTvwB���͗�f��o�|`��"B<�;�i���~c[�Ec}��2/���qo7����;����N���KV�XA���`,�W�^Mh���nVҬ���VZ�ZIL�Nŉ� ΧO�sV��OL6WwQ��	:B%0��+�-�t�䉑��^�p�U���	NVL�`���%T��t��e�j"���)�����=n��E����i����������m��hM��ӔŴ�������)�ۧOP��"���?m�|�[��A�=C��p �������}��	<�'@NMC�I�>_��tsAuh�\U�n]�u�v�O7Mp[�k��O����Ea� d>xNN,���NM��?�R�Ft���L�<{�E�A�������_�o��Ea��{�\�Α��zݼy:����g�>��oڽ��b5�8Ps����P��زn�i��e�S�ۑ�A�D����R�9� ��������}��g���垴��ì��w8}��ڃ{���_R�O�J���md��(@*���+�%��l� d)C�W��rU�`�"�����֭����l��1@c�#�h� ��~\m��]U��[�ۻ�Ӯ�u5n�# ���Kh�־N W4͸�,|��'����~%��cڐ>�е�S�k���t��D��-�~7~R���]�K�K9b�6�Z�U:ӏ��yD�Z��a�8\�K�
t5�T�~��v�J�h,ՖC��0tgsDHy�܍ٙi�v&���[>[�=Ap혅�<X	���ZX�mʇb	�'�}�d>��E'rn�tr�.��}�S�Ry�j��d�3����e��V<�S�~�,-:P;G߯�^]��Ļޯ~�{l{���/�#q� ���
��|ϣOc7���'���;�����*�[��*�<���V�^ޥ����o�q�T�9�Rq��H�m�[}kޠ�#�~����Z��_�"�F0�j�}�������4��4�����{�:7#�'���E��Z�(��H�� ��ڬ�Lp�,J��ݢP ��U�N}��$��QK(��D
��txwil�~{�z+�uﴸ�=��2�C�S϶�|+���T����e�4��>ul�`�{�����qi�l)G�{_4���מ�0_^�2^�l�ٽ6}��;������|dv+Z���L�@�ܓY��t߱��1�<Z���_����������S�+%�y'��Dҙ�7H>���������;�@e�i:�$�7�S�7�Y'sĵIG(h�z����~{:1���\Xj�-$l� ~G���n�~��~�<z֞ONP&�tԎu�9J.s�o�>��Ẹ������{(j����5�RL.B�Ycj
Z�؊��6�,��B��o�I��� ��"�1��Ί?�P&O -]�����-8y �B��W��S�_����v���vµ��
��.��G*3����mG���\��%��o�*�&\7�(\��u@�V���i�ҷME�V����NӁqj�Z�2�5Ņ�Ev�
x����P�;/�-��~���P��hY-ePw����	���sS9��
���)�����ѐ�vH9赯;mz��a	��䗜���Bu���� �EK��H���(�/�Kgwȹx��t�.bY�����g��i�]\^
�d���:����͇���
���{�y�m�)��'�l�����ev�@e(�Q-���� �+ZnW��D��'�}|.Ƀ G�(ő��{L����$���ɩI��ֽ5�^���Yy���Ȍ;9O�e��a�*�*��7�d�Hw�>����^�C��w�騹�,�:�o�s���	���6-��A�����#O�" �J�>�>y�4�uT��d������P�K�-ӆ]�^>Еj������gک3n��ZĀ&�º��U2�7
Oװ��]�̔�UF�o�s���po�h�.�����沝�W�CE���+ �id�K]=CqV)2�K�j����7��鶧��9I��Re��@�R��|��"g�D\���R�n���z߶��?��W�]g9�g�����*������K��m����d�:�{��r�W��Ȕ6���K� *��R;grz��@���l��=ԣ�kLr-vq�A�p�����\˟�)�R�#��>Q>��k����_w��=}����Mh$�3�=���3q�����b���R��]���.2e_׃��F�ü����� f�0��4�{�o���w2_�����:�Q�<n��hY#w��?�&Cj�����o3�v��㜵�޾u-�~��}޿{�a�Q]_n�^p��'i��4��8�n&椱�>D�qh�v!m�0��&Bum��a�Z���=��N�l;��Y�LG�s�.��M��%:�l�#ib�Z�M�u�4��V�P"�Q
Z���w��;9��#g�àjaξ,���6B8��2�`P-�x�ns��a�%����|f�tfv
�L7T����CZ��_#�+�m�Z�3�kNP[������-P�-g-���#������1��?�/$(dz�[G�Ui��]ML���!I�=������k����!W>�ii TR6��u��P��-!��
~28p�����hq�M�.d�
�}�fo��Z�tpr��3#���S�r� ��g���X�����끮B��(��V�\K;ϝ����[mm��K<J�Fnmp����L�o��������z���?��z��;� R��)A����j�O�h��;⢿��y��r#�r�?�O�ȏy��K}u������}�A�-`�֛V���Ȼ���z��#����<4t�p�] b�N֛�Ua�{�������T��!�.�������[O��m�H_��>���?l�~�9r����� "�R�Z-���r�Nߕ\��d����0GGx����%���[�{�]��
&�47�J�A:$�ˋ�:�Zi����_�_�X���B�;쒉�.��m���
v�AK���*\]E��I�|x���'?j��?i�������3��V܂\G��Zm�nP�I�6��d�\ �޶N�	��uc9�J5g�3�a��UA����A����W|�@� ����5TY���D���p�h�n��jׯ�lԕL~�~��P�A��������h�.���>`��Z׷�B�si�( �;*�Z�Nt%���قʳ}����G:���3pT0�ϵuG�b�5�)e5M�5�T֜�Wn4� !}%�.�2�X�ؤ�9�.'�Ѭ��~{ h���F��.�H��&�׾�Ï�~�q��{﷫�/vOƺwP���u0m��T�Xp��R,�9s�e��~����G�w�{�]�x>���Ȳ�o��+�c��>r�bքG$x���YW����QY+Y�� x&q=J�/_i��a��~�>��#Ҽ���������&�a�3��P�����{Z_@�X[��.A�)���v��J� ��ڦ��8b��h��9(�I�Z}�`?e�	ukR�IW@rê{`G�o߹G�6.]h1#�h���
�5]'yʳ�O��#�B��ԭ����vg�kȾ� n�
W�%��A�����~^���.e����k������?����{y�[��AŮ��g�7��������lR�[��U���7�驜�0W��L�@}�ޮ�VK�+��� �G�ڃ{N�@�>�ڲH�$`�V 8�\�2��u��	ON�Q�S{�p0=
-]��j=�/�g�ΎAQ0�P��w���aá
C\s/��N�n��C���I�2��+ڐBFd!�8�uK�3y��$�~�|?��ڡ(E���Ƥp�U6��^v����Q���\jĽ�����v�|f>F'w☳��t�o����#8���Z�*�ѵ�U�j�A���şR��LZ���TA�sw-����M��fw����,��Ko~'�	zm�:�;k{qq�����hA������O�"h�v	�-7h�vB����4�ގP��l{����f)3���\����9�~��uH��D�g�wI�aG ҁ"����p��Q��O~� ����Ҝ�8fg�y�ιB',mМ���Sh�v�ZU��=����<�Լ�Q�=w���B��t���x�P�m��r75���*p�!h�� �ta�����˔��4�,�9+�Lö(?���G���5
ڬf��8�I�Z/F���n���+\���-��Wx�!D�	褵ev��ٹd������xk��T�>=�,K)�v�u'�W�����77���� 0�'��.]��� �V�>���|����g��;$�%-��Z+{?t����Z�^B�I󜏹�Pm�~�r�2���]P����v���v��;�e^`*(q�jgcZ\�Ɲ�N���h��rZ��,����?�iܚ%�Kf9���|N�s�	'~^t99�~�~"���1�^���\P�кzq4m~^����DY15" ��z:��De]U��DF�s���'[F��) ��������0������C��u�҃W�\�J ֽb:�n���mi������@��#��O9���_�W�H�,'��G(�I����Κ|)B@���u��k�j����O����^X+�����S����fc�� ʇV@ۮ|%��b�E���?��d2�(}���p��#\.+)��՟<E)�L�#���Wy@Ru��5(h�u3�G���>�h�ʤ���Q\����e��T�I�J�%�f���&G��?����\V�A9r���O2W�o r��8aZwA�O=�Wַ�
p3亀ӛ��@]�Q֫�,���9Y�)�� 0{�����#�7oG�.pk}"�Kڊ�t�`��u�ۡ��'?GiC�	j�v$���>�߂�^�=��ן�mƫ�z�-Ӧ^�㏔u7�y����G���8�ovC��3/W<����*HG�JB��F�)[x�6c|%'U�_�h���<ʡ({������Ns}�$��Ŕ̄8�?�O��������G����V'�O�1Tf!r��kJ�F�֣�}�u8��3�/ �FGF�L�5��%�������1��{-�^������SgϪ���Lyg�|��G�����I���h��]CQ���f##݆t�XBK��c~J[�rPPC��IN�8І(cYo�������:|l������#%Hwmg2+��[-���d�0��3�]���?���e����e�:�_t��j6�VV6�v�.��`��s5�=����O{}{~�{ꤒA�j��$ٛ	%ϟN� �F�p=B;���
��)��af���/��U�\�сɉ�9��(�'O�NY�z&'�YA�\9�۱	rd��e��{�j&�h1w8�e�n޼�p������5b)����ǆO�S���$�c5R�~�`������k���H�ə]Y^i�[oY���)(�Q�n���R�F�9;|�:����\��x, �/���}���ş�'O��3�]'�ݾ\�k%u�ݼu?�����{?x/K�	��U}6=�(�����B�������
>�{�����_�[��P:t��]j�;c7��K�z��B�g�D�S��M����N�s�	���Qu�Rw�2.���W��h����l�9s.�P+�|d�!�S+�t~��q��_�����X�T�N��yr�zq���O k5D����Fׯ�O��_砣�8qt��rݹm�i������*zgM�]��ź�<]���O?X�J�KEVF���`����`��ʈÇ�R��c1��)���~�.'��m|�?7;�荌|���4�R��UCw�>vA~�v�|�$������9@U��.wt� H�R+���<��I�0��)-��[g֋>�և�ܞsw���� ]��LZ||��M��I[�_H>�߸믣*�n�cGo�ﮈn��J<Je�G˯Z-U�FP��rm]�C�q��"i�n��ׂ�q�|x�r��9v��D:���T�z���kPqwM��W�%��`��&1�<w��Z����8�?��v�X�*���릱 5Y�d�ʍ@zM�'uC7��'�YM�u����j�ۻ%W)�� ��+�P�Ww�tN�[�;)`��u�Pf�ߺ�ԙ�g�����9���$,�֑~�ӓM7)�vY��q�����}�Yc��B�WyI��\��t?8�]C�����y�Û�t{3.e�}�#�ڡ+��U��$�������2y��]�B�,�����㟖�R>����![�#�	t�)� �&i�$V��h�u	8�m��X9�"�h �
���Y���1��cv5�����h����P6�>���\�RbjYV�����j7�Q1Q� ����`I��r��ھ]���{ֆ�M=I=�U�
������*��zx����ک��S����đ���U�lPf�,w#���K�i�R.Zߔ�v�&a�}&�#���W g��=BD�MK�P���;���T�/�`&)�K��9G�Pӫ K���8�Y�@.�~�ڥ��o������~Ծ����߾��{���o?������>6|�>��?z�{����9�����g�����>$|��w�G��r��=�?������o�]A8�$�%�����X�(��g���5c.yW!ng���ZE���}�8���-<�{+�?e{�.�ƥ۔�������W�1p��w�r����ۜ���q�ڷ*����H��2���v^��u����!g��کUԿ��`����i������H�����I�!�����IW)���Z��Q�;r�@�A7����� q���:������w޻�N�@��� ��d����`'�P�@^w��% �v\v�iҹB�t��{:Њ���$�)�w-R-�
�Ȁ�&�ˇC|���(Nh�{!'M��Zv� ��$�W�d-���N��9����엯\l�/_��I��6f�9E'��ѣv���L�2��x�2���_Q�y�u���k�rU��B�}�����h�������K���	@�kESy�v�<x�P>����
>n_߼���� g/l7
6���������ʝ�
ڙ�K�3{����qs%��K:iq�� �ó�7�<���F$�Q!�D�X����{._j�]]_K'����U0xL��`�N&r��zY���T��7�{�+�	-�Kj<S�Ѝ"K(��YN'�I@Yj�m)�������:<�\'����#�9���/ 2a��U�tuV�mِvGpEY�н��ZL�-��w����Io!_.^><��3�A*Z����<]F��|�ܤ�45HyP�9x9��GO�*"�
�`D��E@�E��S�:W��x�5.8o;���[h����(��*	�L��^��xy��*"�-Ƿ�oܖ�]�^��: Q��:T�vٺ���r����+�|��NNffb������P;{�t���~��w��� W+���.u�;JRm栖a���W�ӊ�P�43��.X>6P?y4��U����Kx���L��~��"�Ð	{��G�i�ۀ�5@ ��6��}�� e=~"�����ёU���1e�o��V)@��Ll'&��]#E�䏎��QN�����k}ԏWN��$h��;>��HԅxB�,WvP)Wv��"*�jqWdS�G���'�U�'i��oo/�\��\�ۥ�hW�H�09j�+f�?Ea��H3���K�:퐄I�8���;S�ԩ�!����m6M�e��Ѝ{��-�)��Mr$��/�
�{kud�{9bY\�]�[�/qs϶/U~	:�d�>����5�1x�q]��?�F�D�׶�һ��w� G��������������#�f����֏%:Ѥ D�� �B�Ȉ�N!��S$�0A-t_��-��5)?4�����No��?��)����I����R�Qʓ�)Hk��3t� 6��#\�|�]�x�]�p�]�|���, ���E���v W/]hW9_�^���z�6}v�����;��>�U������v�+��L�@�p7������! B�3�6��<�C.�����r2YV�mh�����}"�<���OGh�o����,x�{Z<ϟ�L�\��u,��߉'ܝlh���"a��5@���[�.��g��Cy�k;E�Vu�aJnc�ѽ�'���P��+p��n�)�,���{��ϟ���rEZg�sM�lN r����0U/��G�J��Y��o��[o_���:0�������=/�;g�ꟆB�v���rF�k7_�v��Q�Q0:�C��ɑ�v��:Ʒ�kYG���`�<͘뾁+���*��
ZU���:ۇ�Lg�UR���Y:�9�a���?�ڣ��c��(������Ν;�KuȾ@9 �O��IG�3���B[}�=~B��ԥ��k�=p����Ew�{6�\S�I��3�ujr}bGb�:-�]��\���5N��Tfء���Kj��w`��]i_s+�R�-�K=\�r)�(�����`�#G�ƽ��C��s=v���n76_X�˯�K�/?���琧�����{>=N��Ϸ��тy�:*w׹ԏMK��j��nWIe�jx��Y���k*�����6��r����l�B�u�,����[l�ኝ���������^:��(Z�۷���<|!mD�l��w2��K���3�n׭��t�����
y�{]��޾k�~�v��λ��x:�e �3:��E:Z�ʑ+-qZN�^Y�q��nd��r���G������%Ȟ>O[:w�����/����9J���܅ȢAs<{>!؀��f���F�÷��T�b?D�2m'7��ߪp8R���+W/S7e��d-�/�������[��@Ty�.]��P��Dɻw��Z���|�D.���?.�O�B�غ�V���Vc��ۦ���t_<C;F[�ej �V%�=�^Z���\.�ftqP�G�:r����G�Ϸ�l�˝[�;,���� ���(:Z�d���]ũw�QɁ4<�χ����_�c��>~N��c}�E��x�;Z(��ӧY�O�9c��_���W�\�<PQ��P�3m-��;�����3������\#ܝFm'U�����Q51�e ��ף��,�T-k�eFe@?U���x
C��v���vں+��u���0zu�E��O��s5��Z����H��g$��@T�!�%!e��ɷ�T�E��A����P��www�Qz���V�)��d(Sl|�;�q��h ���r�b9��s-�b]oȍ�g�9�-CO&{-�ᡘ����r��-&�O;�/�hVF�*�G@p�ţ����a�s�-&��ݾY٬5Z%��܌���q��NC�ʇ��[�Ǿp���ܺl��=�@�`d�7]GM���LtD� �g�d��Y���^P<D�,}dGR�
�ku�-��k�>�N���f�|�`���>��۸�N����*g]2<�@���H��0�9������{�n��w���ܹ�u�Z �:$e��ڽ���V��]�0�Ttg�ډhEu[̳gk3�u���8g5q�Lt�0�G�hpK���^�`�,S��2�<�-t2�.
�}в6��C���q�4�Ut���Ե�~�	~���A��m�6^GF�B��v��% �:v��|w�~��O�8;z6tT��;��@h�u!t��tMG�l�y<�/�::�갤�)2����߀ũ��������Flp�U-po��UF蔴�*H�v�
A���|��M�]��qI��,���m;�Z�&V1�!|l����[c�t�Q�-�?�'-BT�*F�c��İZnh��]����
7����F๟6�Ш�G���6���=�����q����uc�Cߴ�m@�k�>����	XO�<	�nw��Gp䜁n�AN��%amւ|����y�N��v��F;B'w��^��dRn���$�`	\�_W-��u-x*;Z�tUq)�Ǐ'���ɩ�.�_8h��/��%�	D'���ɗ��(H[�]d^� o �����
G'���Թl>p���NO/�;���`�\bI����'�:D�b1�B�D\��*s�ȫ�[��-xQˠk�ꓨ��u������̥����ժ�ڨ�Hwb�D�()���ہ X����wޢ} @��]�x���.q�mR��*��@D<�އ��v��	ۻ�wn=���Z�c��n�B�O�E� �	�U]��w�3(	�u���
0\����-��ۧ4�'�Ia�B�-O�6�
�J�����Cs�2���z��i�^̷m���e�zтYʧ#8�,�4�ܞ���^�|a���e���V�wXSYp%��v���N��M��`�7��wR+<E�$�w ��?,�9�+?�
��rh~jJ++�|rd`(mT7�����`w=�/���J��' �9�Xm���,��_
lٮ���ue��=᳧O���A��U�tI��a;�;Z@��V%�z<3���L����2�>Yc�ʁmCѝKu�qI��lౚ|?��N4�<օ�����>xB��t4u�YA%����w�_�{��(�t?DŪ�϶��m��r)]�kyD�!��!s�B]Q^�tm����I�X���?:�N�%�7�k�b��>�Zw5P[���>�M�gN��Q�6�LrB��ۿ*�\_ؼ	Z]1�2���^��V�����
��N�Y>%1��4� �]��4�|� �|���;��:�_��N�yD)I�.�%���pY�Y��!v2���Q�-�A�3Z�O��}��
�r���_�������Z�a0Ci4�n�#O�e������.�����)���G<���T����|~[H+�N=���T_UHҐ0H�|*�3�!|��[K�����{6~�Z�d�.��j|�;�g�i�t'���=YZ��1��L�9��R��.�����
Iw|l#G�%Ѫ@�A��ZM�It"�A���A���V��� ����̰��)h�o���eq���]��7;���?�k�ʹ)�S5���R6�bL����B��ݫ�j?���Ȯs{j��`Ca98���	�kҪM\�^���\�|��P����dZ�t�cd��bt ���@*�W�^B�)�yҵ	g��a����y��- C@j�ldoI�+L�N僭�3L'u(���qI��St2���Ч�����`՚�ց��Kth��V{��w����Y���c����#-;?y�L:����2�������C�;�I��gδs����.�7=��F�Czfך���X*�'ڥ�Wn��*XXYy�� (*p�ߢJ��q�Nh�t��A�Բl���v�  tU��&`_p"o���;QQ��=�_J��[��ڤo�[UgR��mK���m?x��� S!����:�v�ݿ�8�[w���J0p��8�c�=�����ю󀊳QVͼy�|>�aC�>��?z�N�vڟ=�wt�n�+�9��ӹ��7�Q�@`�4�����: �<ʷt���ʏ�^��V��bv�r���t������y��e=L~�ڄ�P��,�?h8u�	c�zt
�Ɖ�g���Sɫ����F����n\���z�"���1���<s�}���׀�Օ5����h�k����r�l�P>e��Y>��8>q�Ɛ���������o��gU�Q��7�^Q��; Pt3����2]�	�,�V���~�w�Je�tx��J�͑�������F{[K=q����������щ�Q#s�.%-�i����>|t�i�Zݴ\޿����;BY΢�\`�� 蚝]EM���qÙ'���8��Ѳ���+�,"��*���*��c�t)�q �-.nA�%�����nP>����*�:��c��Q{��
|�Nm3�y��5ʩq��E&g�R�2i��Q�;<�Ri(/M{�tf�<��0���d������.�O���v�z=�
 ��}�]�6(/�̕Q'Ojp8�FYf�n{����vw4�@�a_C��vR��G��A� W9�����y�����! JB�5�@,�H�@�&�es�SȻ��Q�[��D�X��0B��mn��QN�k����d�O�mF��[�If�����̚��+��+�m��-�gϜlW�BY�
ӧ�ҍ;e�J�����uڈ� 'V��m��t�s�'��h���9���Xi}��{�7�d*�T:r@�^�2�aG��W�rϣ���n�{��rK~�蠡C>����u׾=L��R�Uy�:���&?F]LR�w���v���wG8Q��!{Va%���* �f�#se�O����������ّD���N��uʳ�{�uC�k����L�>��}}!���ㇸ���B[0[�q$�eP��3)l�t��T�m��h�sY�+!|SK�m��
t暆߇�]4��?s�=B�Sc'����-W�D�Y����+�D�bz.����˫ۀ���$�օ��jfy�����g̪��L��iá�
��.�E��cS���K�����Q�ѡ��.���m��y�`88@=� <�,	��x�|ېv�H�a�z����=y:��C�v��Th�@���m������Ľ��9��5~C�Bi��IOX���n	�@tH;���P���)�KeV4�[Z;��э��;�NP�V@�(��� ��}v�B'5��JRVȈe�ɒ>������R;}.Wލ�R���j�ti!'e	�����s���9�T���籔�' p򊝎��m�:�iU�F"K�j[�I��X?��XV��ϝ���A� �A�5�z6N��f�����ɹt�s[a�ϥ������g���'� ���_�e�E޷���d�
�Vz'A�'x�
��zn�룇����:���a{�N�9|����"KtE�����拴�:t����������>�L@ mwy^�֢SV�3-�/�k0���M�7�M�6�Wy�牰�<��reZ1̓��-k��f�'��?�>�\��t�8s�Lܑ���^'�-/�D^�*J'<�/�+:���4t~�d�| �]�S���˫��g3O�[�ڹ�<u�����?����D�ƉUT��m��b�����PrsF���Uˬ��n��$W�g���o������s�(t�n�z���H�B����3�'��3��_/�[mY�;���bF��)�(4�<ۉ����w�2؉g*d*����c*w�H{g��B�﷖Sݿʵ���#��n�ew�t�A��X��#�y-�ƪ�Y��n����f��}�rж
!#ۢ��Ie� �r�5�����%��P�������.�ԍ�8+� ��k����^��6�!^qe G/��+��,���9��o.���Nk�9;����܋�V[yn7x���/�?�o������u�u@L�j�GV]�ƍ[Π�n�����Jh�&ا����U����/s�f��W��<��k�W��c�&��
V�sC��� ��:p��@����5��X㵯�5�^����-�A ���uzw�-�Ƀg�d�BN�����<�7�~Σ�����%>��M�\�+���k�����v�A���J�[�Y�e0J7��R�֥�K���#n2ጾ�������$�d�w���Αw$?�����߱���'����/(�Qxϑ�)�a�0=Sͮ8O�ݣ[ﺃ���.���|���:�:�Eh`����;����;�_��[/�r��GMf4+d��_βbj�O�`PIZ�^*��c�:kTp�p������v�.�p��VÿKn��o�������^{�[����1���>_]��痴\4��{�'n����V��7�%�
w°Um}�q����� �Rb����f�W�Ӳ ;뼶�t���~[@ܵC�H��t��ȇ��F�������xfV�m������ݧ�\�� �-4J��Chwj�
RAm�E�����<�X��r&B�����8�(�E����>onb��QmH�*#}�bC��_7����0�C��R_�t�����T4RBiC��#��C�����E�\ŗ�ƫ��ȱ!:���O����) ףv�{��Y:*'�im�T������X ']VVP h3����{jj!���-+�P���5/������ڃI:�g�.4�}�=� �\p�����QA�@XAW����v�(� Zӟ��lϜ`��e�y���s��m����.>|��-���%Z�k�|���y���]��<�^1�n��.RϟN%o�I��t(�Ӄ���>��Ct�[�
�@��� ��j���y��ҥF��}!4� �	�vVa(���Cv��l(�C�n�y�d��i��bۤ�:r%�V�&�漏_FVM@�{ �/��K�<$����6:V��qxs���D�(��K+1�G�y������ͭ���C�0�|9)p~��T.�by[_ӏ�p���'�P�Z]_�E� &�8�/�^h�LH޶�?�rSwʙ�r�4Nd%
�~��I8�k��!ރo�������֑a�Ӯc꤫Įm�goY'-����o�g%�����ē�7�}����[�[.�����+A��h�!CE�!��J2��ڪ�#��J�W�[Di"(MO�<K���ĲT�mG�"��v�J,���|����[EH����������}�n�ʙ[īl
X5f8*���נ�S~���"��*��Z�G��c��'���8�`+m��]� 6j[�[�U�����h6Iy#7�{F1�^�'|R�!y���H�7���Ԇ	��h�v�[�5�j��胇��~�>�����xJ?�>�_`�?Z[d|�(��ٵє�Q���S���(�C(R�݂�lpk|P'�X��lt��bn!����l��xOL��xY�g��NݿBSf�� ��^�����5"�۫�[�� �<8�GX�k��U��H���ɔ�v���.����[n�H�P,4�[�����hh���.�Ѯ�i��q�����~����U֔ڈ/󯣉�6؀�[_V	)c��td�t �~C�rK8�
n�*fe:	n�����|���L�K��R`G��F�+��g0�R�
�E�s�K�����3o��{�\�e;')����k:�D�*�[N���ͥ�V��3�Cc��*��� �b���ſX	!��C��O��_wLmfw�1���={?�$&�]�L����tkO�!vmͅ鳫ٚ`��H]��6;����t��"w���Ŗ)�+��?��a3�T�/�e���\�ۥJ�QP�-�]'�0g�1T���� �]b\P�� ������gU��u*.G18y���KN2�����L��&����5 �t����j���c|����ݵ�e��}�_�~q��������� ͡�c�%���F0٨�R����$}�VV��V�E݆���I�Z��|�Oq�Uw����6,h�?���̇Co�ղ�@x����O\�Q�Ɖ3��MaRN���%�N�/���ڻ��\��ƍ3�}0�g;ɦ[���)���V�t�0����R{���\������#�al
g�Y�����;T���K�\�t��:]��<\�yup�n=�StRvPZ��,]C؉p��@;@��۲��7����Qf���ٰS�噶��M�S�����/�=��*O,��OB���v��rU����ȶK��m:��p��ԓ4ӝD���l���L��>z�02�V�����v,~஄���6~
`��W^��PW�Qt �0�~}���'����{���_p�*�� Np��������;��v�n.�-��ʊ�9�i�лÌ�Ug-أCqKpM�3g��ؘK�d��ٍ�i��TW���Pyb[9w�T�*W<p)2'�9�ffj�͢H����9�(JZX�k*������,Y�vC+זQ�Y뎶Ж��y������KG�
��)��n֛����ġ~�����D6H�l�3�v�ӹ�(U�+��/\�w��ptEPI;��]l�#���&�e ~�������$L'��848Ԯ^�W����sn��ߨ;��щʦm�e��Oy��Z[*�����uG�G㱿�Δ)+���s;	o��slC�r�e4�5�|���<|�����>�_j���+[@V6�X�����[ �W(F�����.����/ho{�� �`�}���C��MF�Z�Ζ�Q�a�=�eэ��k����z��J;�-ВN�sk�I����$eu°�Gu�Yy�e��^�>7�H=��/ȿ]�4�|�� �Æo٪�
W�?z����0��E@���84��Y^16(�7�_� �7�����Εx�Μn�s�]�͜�����+��F+aYucT�;2 �wn�S���t�E�]C�;td�A��ltT��U�Y��u������w����bs�m�L���}��ճ�G?���ɟ�q�v�2�`l��_�|_Mtx�J�G��Xn�!x��.k�Φ�6������S���MI��Ռ�Jh�R^��Д��^�\�ĳ��ST(�[(�y/�u �`����N]x���+�"X�����M0+L!Ϗ���#���	h;Λ�}W���&��Z����v^Q-�N>�=v���������tX����,S`�m����K�$�,�#HL� ,8�=+�$�G|BDOj�Z��8�#4^#��������^*��\�ù*����/�� ������gV}�� 㫅Ʀ��.!6�.���8mL ���v0C5h��a9h~<�4�{�Ȝ�9�݉\E_�d�4�O��P���e�
�GM�����ﰟ�	5r��
v����Op�è�>$TW������XP�[ �}��!@� ?���(7�UR�����+��q�[�����&��Պ+O�'k-ï������smZ���n���}U��iR�wV�M;���d�(��u �O�]�!�)qZ��Y?N-�.$pҗW'}��`��ix�P,BVw̾��nxd(��N�Tٳ�Zv&��}�^���+ˤ,��Y��� ���̓nֻ�
:�Z��M<�j����u��[�
-��va�'Ul5z6��a:�-�+�>��n��-F�~�g����x<��j�򶫶�na۱�-Ya����6H�ܐO�>����Ln��xi����h��!׊\�w¤��I8�7�����I� Od��Ϻݎ&l��Й�.��v�.I��0�S��̞���Ԑ���K����Z�Q�>
֣`Pe���ఓ�ہ�!~wtt82��T�ϕe@�< cz����Qv�6K&���>x���<u�7�|��.�҇ORC�Z��6�U[Zrk^@�ȩ���u�@���6eS6:4��4��+�]RK�7A�ҾjŇ���E�6�(�g[��G݈o�K�FG����!`�����c��U޷�_���̏+m���}��i@����>{����yQawƿ��圤���u>��̿��ȣ�,OHy�K�EA�&�,��k����E�lJ)UTƮ.�7������U��k�'�
�%��?��oo�Xl����K ]�0�t��H�p�P��~�� ��]�,��H��'2�s\�����b���ml[`K��g�*�*�w�INk��6�T���+q�s�2(O��.�6�4ً��=�7��[eJ������i[�����;���֕i�Q���~�<x�]�4�97��!���^��H{���ٱ6�\��
��6>��֡ Ց�e��u��#P��U��H�~�.�Fs�v��{�$} ���[`���n,�M�����v����C������i�U���*n�=��]p��6"�=u�\�n�_ne� \�I��S��)��?����I��y���T�Q2�� �������g�N��fī��oۙ|Y!�C��Ё[�L}n�Q�`���[����1?��?�?���t�s��]��٨������ay����m��A�����Âʘ
��v�aL����DZ���eG���!��#�o�,�Q����Ep�O>�m�o��¼.�h3NE"T���6=A��������
a�i͋+���`"��7�2Iu�q� ?�W�m�-?bH�u6�>��"�:�۹�ND��˔ٲ���f*/
�	�e��"ۙ�ĉ`"B����8��_w�d�4��+´~a�}'ޯz�'q"t�Z�Z���b�w�z뱯�ZR̲H_�6�Ѻ�N(��G�����U:�c��� [�]���[��0����$�ȗ�J��K��C �-�IH�L���=A-�Q)�3����3A������X����٣�x5	��^��A�A?@wm[B�-�1��ֆ����0�	A���?{�w]�[:i��t�u��1W�8�;˩E�e��%hcM������3 V���%��i��Ey:�Ҿ:Zx.��9<��h �պ5$�m]3غ5~����6�0���\�5� �*�V�F��>�G���oIO�-��]�%�"vh�P���ɗp�,��e��Xqߕ���9yU�}���ۡ�����v_�^��gZv�P深�� V��6 �s(�+k'+�k���?��MGã�<�����A]�$ض�'���-��m;�6����U�ÿ��,pG���.i���Ҏ�r�Cw'�:��jS^�S/h��U�ey@�%(�;��m�2H7y�hL�@ਃ���憸v�p71V��g�C��w� �8�UQ���U"]:M��;�ѵ�mYۘ�,��s�:�}&�B��K��]!?�ٲx� �ܓ���`>e���Gޕ��W�����r0BG�y�k�V'�Bx<���!�=G�W�>�!&��r%rФ�4����R�򬲂z��)����CBf̷@*e���c��{H�ޯ�m��e4�rT���(�a����n*�,J��Qy^��H�-S�[�i�җWˈ��Nn�"܃F�-��vT�� �JԒ�*{�k#���SGۍ��ڹ3�ڱ����)_�c�)��mO�Z[Y�5n�=~:ٞ:A���|p��R@p+��}�?�B�h�{�|�<���N��v��ڟ����W/B#hx�?�P����1��t���0J����Y'�j���f ��XOD@̇�9){�Y��m��R��V�w��'���2�B�p_ߍ�O�g��$��Hr�k_�Eے2�x5:�&�uc�������R�q��B�'2A�r���:�������?��uw�sd����� (x*Z%��&���]D�e�{U��4-� O�	�;�ם�����3��C�@^`�����{~o<u��iէ0'a�ʰr:�Pp�����p��dV�����X�Q��y�w�ԗ����o��o����?"4~���N״�7�u��B����'�1�t��7��{����+�S�ҏW� Y�g�s���KuZ����OO���!�:־����>�_���p�
P�]"�����E;B��n��vp;Af&ɷ{��u�}�Q�_G���封�l�Y���X� 4Z-��5@f�-B����U���G�/Y�di~���Z�H�Wխ[U��i�a��0 �4j�g���C�` l�zЪn]-���	��~�r��Ddުj?���v�|�����F �Y�UCQ�x�C$(�E��� ^��νGu�[�+e�xV�����J'$x��JJ�9����JG��J����ぢ��Q���T�W,��q:!:`�#��Q�����@Н9�ҠZ�*�u�I9i�S��HQ"lg7�(���#^	v1ߚV䉃 �)�	�ş�(:�8�P^�r׷\��6�XJ4�`,ܬ@���x�G�t��1��-9�;£�0�:M�9Cipb���I��t��P��(Ԗ�M2�*�=�����xc�t����l%~�z����h�H�nE��T�إ�!�6& dh�-¥�N�(*�>�M���t����th�i�@�-J���L�<P:jk(<�#u�J�'T>���(m�ug��C����?�_="�q�����|��<<�ܴO��۝��&���GyאϔM��hʒ><�?n��z�ˁ��;�.�����"0���]�QFp�%}+���j<S���?�8d�q 1.ԭhR���H[`	�E��f�۸KÀ���&)D��(��>�!3r������Q.��nz�\N��8ʸ��]��6J<j���`JL#�Z��Vz�i�(x08�oX?��_�G���\$���%Z��¡ I�A�_�H���+��n���ܲ-��⸕ۑ�^+��8z�\�A���"�N5��l{�W7v�i�H��мP�qM�0QTF�m��ܙ����Lh���{i��UxL�_}�Q����*�vN���V��f���1���!�Q��V�<U�������ׁ���L�T~lS�<)\���g�+@~.��A�ׁAш��#���!MR~�p���+�!�� �|E7�b"���ٖ�G|�U&�������}Rn�����$V�Z�O����ow�9��)e��0J���7�=#Y7�9J�_2��(~&&�҈�!M7"��[���
�2�м�x֏w5+I0�S"���+e�<��j4���F�W��ʏ�]7D A�N�9�8q.����P6�G Y�<D��|�N�2�g�R��o[~<7�+�Б�.y��!�kfTכ(�Ѐr�x�.1V`����T<�w��F)t��)e��&?��x*�$@��Y��Ψ��i���T*3��МO��"�R"��*�-��;��%�彞Vn�3�JR��IS8X��  e���	k��\&�A���k��rb�8>9�3��~^f{.5���ͬ���(����lb����iy`��%N�s8�C�p��ej��`����k/�}��rr��|�41�0u�UV��t�"f����4�f�7[�K<фQ�7�s�:�k�q��H.����#hU�%�)~=��'�u��a�q�ەx��BQ�]�̉��	|�Ò�]�� ����i��dx�������	�\g�'�'�&J&���#8� hJ��>���ɼ+����傃ZН��lU���s;��Hu_�M��6�%�����(;�_*����#M�⑎�D����A�P��6沠����d��B����ZEٙ�f�� ~$&�2�t��!�K�F�ekP=.���ʪ4�k�	�c�^��B�(m��r[��=�X����D~���r����By�O~��h�6�[��r�0r#$Ϧ��H�)q��Kr�r�G�5���q |��B�!�Y�R�TN7y�E����U��u�l��D��H������/(e�®�̟��<������gV��C����oH$�����AF���gP�j��I���`��3�b��L.+fL���Ζ40Е�Ǹ��{n���%p�3D�1���]m�z��N���g��x���&h�,Q4��<G�^�R���Ko�Rw�����Ը?,��Ҟb���2+K�9>�ͪ��������G���#[��M�w�
�[~$�w�K�W�q|���@}��y?���!��/��`���d۱�����$����?<�v��,s��[x�GMqo�w������=NT��+0���
#p16�)��nx`�P,3�ֻ�
��]�fT��{	���M!h!�=KGCuZ�V!����+ƛ�m�1�Sc&� �n�(ij`Ң�	���4�+h]�8ЩQ(`*�G7@��@P�ؗ�^Pl�H9�mw�1q�*+���2{�;�� zWx�09-C~����'��sq%"��.��p�\�<�.ë�%l�CG�I^r}�~cpBZ��:��1D�H��;f�P.�e��t��-t���iPt.��QZFA6 �͋�i��P�3���(�DC˼��'\��N��C.Eh+U�ი�.�Uvf��3Ⴗ������1xZ�i�Ta���&�P��aY%Ey�Z�^�o3?u'�L�,_�#a@?�I��4�{��<�-Ŏ���q�E�2`p'�ʓ�$�=���J��A8»Z�
��L���x��A�s������.�~�l�F���b���u?�݊��0ҡ��@ی�*���Q���J��e�	^Z�+7U ��&l��0�s9��:�^��u�f�(b̄S�P����?II���:A�f���4�%��
����G�@�ۺ̫���K�CU��0�?���L���hP@��t�qȐ� ?�Ke����A7��l�ب����)������mEr��l��ϙ����%�\n����_xp�����q��sys�����d" .ɓ7�_}�a�>�ѻ�eqy���Tpf��i��8g�'�(��Ó�y�I<�e�ҍp�*���e��L�(�B����uyDX)�!u2���ew���s̴+��1E2`�	C����]�M�g��F��f+9�rS.)�B��-g,:��K����-c��>(m^iʦL����"?��7B�j�:��hN�K��D�'�a�-OV��ӣ좁��ɖ����MRn�@˘�[_��(��]�^Q�H���r����>(�\����L�G\EȬ~��e���������8��L���!���l�7�h��9�����3��?�ȗ�p�{]����IO`P��CoS�b�>C2Ye��8�1dڸ���_c<��Ҩ�8FM��T��.�*υ`n�ƉF�� ƊU�h�VHiߢ},�"\��Y���k5T�����Kn��-�PفC��3�"(�t"��tYX��x�:{diE�e�@)"*W���3w�:L	o�F����L�M������t�{�`��u�.uR��z���\v��a��h�A�h$Э�q=�_P-�'�Z��A��>P������ȃV𲱔-/])}��i��f��)0�{zCY�g	�����U#�2��X�7)3yo3D���b�t`��,0u���NB~���������Ci�%��i���e�*�aBa` Í	|v���/
G��&f�20���P�cf�5.W3j�4�z��yI��|�8�ڠ���H˼��Bd���&��hŅ��1���@�P�X�^�%hhe��W��P(��E�pN=��ΊEP?���Fo���Q�Y�)�p�'��N��q���7���#߰����<�!N���T�Y�+$���/~x(7�2�Ћ��7ˀ�MD�,Z� % +����Y���Jk�� ���e�@�E	��+|L��&�V��)�-�<�#\E��%*T?�3ݳ]ѷ�e�Q;=�o�g>]�A��Ts��z�U3ťNH~@'���W�C��s���YohL�����s�58�f)��
'peP���e�q�/<�y���O��;񼭂�0��Vn]G�Ǡt2���:70 }���_u��^%gLg�ā�Y? ���C|���=�:�@3�l;E�í��jx*Ŭ.�n����M{>��$�d�yUu�?2[ȶo�C�0aW�7Rjg+��ګ͊I|6�mM�Ҁr�-C�� >x���&����S���cǋ��.a��Xn�����	���M駁�9���2��w����vĉW��R�#Zy��Sдr�[��Oq����*�пLng�E���2�3@q��
D�)�prsAi���>�v�jT� ����L�XQT��	�S5ړ<���N�X�����7�\�>�8�N�jd`�0����Wj,�))��y�qx�aW��P�w
 G/�FwM�Hz�8I�5��齦��K ���S�\ׂ?��F���KſR��K���ޔ�R�.��ƒ�n����H�,Pꗊ���p*�6� �2��� Z}��<�;tr�bH?�����? �ĳ�qS�#��s$� ��x��7��G9�p�.,W11x�[�@U��D���N������[�G�i9���Kg$����Aee��V�ŭ�Y��J��+�����_�,kL&ӑ�T�ѩ�D��`�]���)��i���ʠ�҈�<�l�(�<#���,���W��BP�8���eG)��.e���2�����3���	\4ozu���|_%l:D���YqĶ�A=��6�B3V��N��TOI
��<j�y�_�1��AP���L�R(�d��e� n�J�ڀ<�U=s���l�[�(>|́��E�C0���O	�V�+���Q��<�<�@��נrZ>5�rus��C�\��Yi6�/�*�;�
9x1�4�6.��_ig>�@9�l�B<���d>"�mѡtZ̼�x��\r�MgA�au ?hG��fE�:��������7]���yp[h-��,��^q����
�x���; ��f^��n@�5h�OO�[\��i������}��C�_�%�p��OD:po�ce��h�\3��g����2#V�b�H؀Wf�*SP"���#�pE�E6	ǑQ�DC��L���E}��}�4���������|�ErAr��y;
<�<��`L�C�P�ȝ�eP�P��}���}�:;�f$�D�j�#������o)&j\6E����0_��#{�K�r��K\h!h ���.�Ë<�t�\��'Ju�����?oJ8ھmx4����������,t�O^5��0�(�z�@G&7"�$#a�4�m�OF8�}�|�w�Ya�c�x���(���39�D�kB9b���������reh������&e�M�r� ��t"��gHUYNv�ʠ��g!Rע̺C\	j�*p���1�ցM��7 ����{�TFN�r7+Wc�D��LC�t3a�!0��B/(�{���@�P�T��m��)��J3^a��(`��g~a�.#AQd�2�m,��Wy(\�-��D�v@|f���>�N�j�p��ux��ͳr�pW݈�t�l�[5ԙ"���&����م����P�Q��=��O�<�+�O(��&�.��� ~�(�,g4(m�Ԑ���[ �c�4 h�nSy3k�x��3ffq�24�?���RQ�*�𱯕� |��@ҳi�l�#�9��!�V�삯09\#����%X�&��y�_P)ȸ���[�@�4����l�n��2؁�< ��¾r�I���p/
��Jn��3q���q\�me<I'+��U���)wb:oP�H��ʃ/h�r;���3�U_M��z�NJ=f"�c,��b��i�c����q2��@��kN!�,�N�V�J�c�w���(ubP(����\��*|�1#k���в��M��Gh�@��vS��+$(u��4�%�!rt|7p�|Ң�d���N|Vy�����.@��Č��=Ҧ &diC�����-O��a��w�rĭ�X�q>�����O��&ܑ11����v��Ʈ���[gӽ��i~~�w>wu�e��N�{�}����w��ϗGn�ᚸ�ɩ�ԞpC��k'rSX��r��I�8qKir������O���I��iRJn_o�bk��ũjW8�=d�l���"aTV��#b�U�WXˎRgd�t�R�׬�[V"�Y��ų�gp;���M	�,�v>�ar�%a�l�f�? �Pó��wU�/{���Ŵ�����-���PY�T�('��4f��	�u�b� e��Y���2S�7�Xցw�s<��4��ؔ� ~.<���4"����u�����r���)�����O�r1},Q`w:�5jSGՆ��ΕM\9ý��1��@g����8<�)��iH�/�[#�2A�(��YC���V�Ee�ϸ5�=b���lQ���t�b#.���	*[��0���p.�q��@g��U L~.®2��̅"�����x�)��;ڲ�v(�,���zw܈��;�'��)��#�mP&Cq�f����ee��	:���4��)�y��u��.��[ԻQ�\��(�g �q��T��+a�K�`U�����2��T�J#�F:
hwh�+x�3�(�
g���ұ�f�q0��BG'�qg��3%�����F�t�s �����0^��7��3�r1(��JיȔ�m:���t�"����r9V�K��Ζg9�>V�ԅ�v+�1q�?�"� ����߳w�N�s�1�Co$G:,�N�F �E��<
�9m9o�-��d(��r4���$&7�o"3��~��e�PJ�iM(���<��gi����4�����s���zM\��D����϶ ��������S��ЧئWV C^��3e̢�U��M�g��s�8U>9����߶�C�;���UF��O��3[@�Badj���G�F:���p����0n���D~�i�~�/����Z�⃳sw^�n�J���n<�?���L<�\Ц?�K���A<@arXe*�z���p2Η #@ܿx�w�����8R��!�_l|.���x�Ѓ��^�]@�d����T��m�NS�c����t��������+����c��tK' H��?����V���K�R^Ok�%���� mnm���մ���[�)���Iw��K�s�ixhD�D��c�K���rG=O.x3�W�|%mzzB��b�J������Ž�(��K�?��w���ށ�ώ��R��x8G=�r�v�"�?�b�*�����;�Mf�{�R�9���f������ و�>�p������O�\6hK��L\��~P�[+U&V4A�7\���K�=N;�H���-H����0����j#��P�S�8���"���a��Q
���ns������3u����N/�@�ʱZ���,� ���I��0f_���@W�s����~��b�A1�"��8�8��`��=4�l���:_����`8���3S� LCX�N%�qtM�W�ߔz{;�^o�0�|��� �T�K>7���?�%�ʿ=���-s϶;}�<���㄂ŵEn<b�3���6�Q��s��+��(5�`�L^V^d[�9�:�F/8EȠ�8����+B��%X�em/�ڐ�:�L{��ҹ(��V��#l�;B���B���I�Ji����i�%��X	ƒ710�O>xc��s�`���Gfe�q��V��^eP�8ӹ�9�d��m��e�߂E��*_Z:f��h��ȁuD2
K'�gyHÝ9eÙ@�]�$'�Yђ�4������{�mZ
�s��p����o�d'�6R/�s��P�t�Dtd����.^%y�.�j!�FzP�Ȉ�<Cb��{Y��/�|;�^���-�t��4V����/� �d�e^�<����<�<�#��
IV��S��e��D2>>��`���2C���~U<�ɉ����H<�c\�5�c�x�l�ď?�t[90&�V���@tܦ�ҏz����$������d�+�Mx�E<�}�W�`��:܉��/:��
G쒖�
W�
�?ݗ�@WE	<I'��P�.�L�Y��v�������3!\�?x�|�8r��+.�a=��2}X��SJ7�#x�㑘�O~��U4$R�HCvC�4ڄ5�+m�c=2y5B����n%@`yz.�L�dsU_??7�?���,̦��Q�"��C��V>�B{����7�p����@���P�gp��S���J�=��H�]>�.�+�ž]��7??�>�����q�A���v|<E��.���fҏ��v4	�4+����(����?�ꭔq�Z���-�v!�������#e�-�����r��h�+��1h�H�������jٸ�6h�J��6TdB�CKE'�����8,��F(���;�}�Nx��R�Q`���S����j����������g/�ғ����枯$�
�����̟�3��?�F�	5`�O�A�^)[(m�|}����-eV8�������wu��؜8�ie�]�I�w��$��	�"R3Ha
^��؀�c����Ejk�N�:Ka���H��C������ǣ#� ��3b�5�S��<�?īz�O�p�$�imu+=��yZ_��HJI�ho�R����8����d3{tf"6��-o��Ω�q���p\[���5"��J̠���;Y�ŋ��&3��e���3�����I�Z��U8=��w�4�'�Ѡy�Q:B�䔏i�/L���p�	�L��&B��
�%�{S�PP��Ct�(���Gy2�4r,.�^MFx4<�$���R��,w�^��HW6ɸӧ�� �� ���ً놥tE���k})�����t:6���1��^I.����I3x�E�=��x(ǲ��xP}�j�����,q��s�9�R�{��(ܝVt�}K��6<M�h��+� h7����`X�-���I���H�����5T&�$`�.��Ao:���p�����6����3����G��p�"��pC.@?+rJ3���|r]�B:�Փ^Ƀ����pr�1�"|�C��8��)7%}D����Eہ'�U<��F ���y�&�r���r���'��'�Ya��<�F�Ie+J?�No��c�b=L��������#�������S����� ��4Qn=�!W<�g�E1�QiJ^X�s�� !�c��3�����N�稳��T\�]��C��@����Xi	�8��DW�;�!&,*�G���Q�~�Nz����'�($Vw���!��	�)�=H3'#����ɗ���΅����k�)i���2�N��!�����1���ԨO���1����̤+��RnC>�y��|�D��F�i>��
��ǨS�G�ĵ?~60���3����(#�+��\��wLI�'h*yzŗOU���̧O>~���7�Hs3��x[[YO�?�}������g�|� _�c�wp��6�Ddt\�m)K�o�g	����1��_��rٗ�ңǏӧ��,��������Z���I��,�z��j5>���Y8�e���A�8��=���Ϧ������?�o�����]J�;�R�F�g7`s;����ۿICc�ix\z�ܪ�;E����G��Uf5D�̭
���.��{��*e�|��.^��ep�:v�z}8VD��k�m���O<�^Q_j�^.q."�51#�O�&+��3�ihd$u��8M>���U��N�Yﮞ���×;�|�o˿��/~��̭ķ���Q,�Y%
���@�npWr���ó�3uLN��Q)��BPvG�>�QȘ��!��h���H|����)�l��.�=}��V��"��O��	�xfm;�y������`a~Z#�I+�#i|l(M ��Gx�ߠ܆5�N��#z��o���q��r�����m1���~S�IX@��ޚ!�+IP^����	�U�0��ܙMw�ۜ�ѱAV��@l|���ö�w��u�y|�7
;�gL�����/y�.���!�R�B�l���aU����wwf��	����n00;޶r�����F�TW:4 �ITW�/�q����'��L��ҸBO)��������t�!<Q q��1�oJ�z_�n�'_>���)��1F�Vx�kM�aT�ȑ��Z�'�VbG<]��h��xC�-�ŝ��Gx�c��t �[Q�;��@8:U��qng�C���-,:\@q�mt�Y:����ܘ�r0��Y[����t�5(�.3WN�
�L�A�p�ɝ�v�"�����T�
�d�ρ���I���CdWx�8��-+L�?�J$�E�Uy(u�H��Pǲ��k��G�{��sx���E`EQi1�Q�拺�F�0��Jt�K�� ���l�(�_A�S8*m�v�����l�z�K�1٘LJ���8:t��?�G� '�s������ؙ�$fk���M\ �����(C�I�I�&?h`�����(I��͞��i� x(���q�N6��Ԑ;����xI`Ў�w�sN�3�؂؛-.Vn�8ʲ�F����_��!l��i�<�^��TG.��qx(,�T��zr�s��� �r��\�H7j��*���gl�b�vk�k���q'����#�G���D��̂��t��]�I�-�O��vr�/:nn��?TVM�=X���]�kfC�j �Wq����L1qu.�w�«��������t��]=�JF�K��P�;ik����u��F�{�d�5��H�n���gn�
LzIʋpb�7V�B1_:�n)ylK��5f����̟f���Y���"�#]�1��)�-m���獶���W���Y�I�_�H��6z�K�(��Z�*za�U����b�)w_�A�3y�����K+�ۻY������ӒE0Rf�@��h���v9���B8+���5�L����f��d��yZJژ�ۡA>u7��q1��b)��|{\�����q=�}&��%p¨��B��y�����ɑ���1Ȭ4�1�?���z�vw��(MJ��}=��=����cnH
6�����������<�8k��鯅�T�f`�Jp1V�vV$�(9Q�b�֪ѕF�����8/�[J*���f�����q��ƥd��Π@�>>:���&��y����x��(P������d(�t"�)��D��3�a̠����ï<߀*l���-�|D� ~A��Xʡ��B����$#gf8��S���BB|���ш�Q B%1���]�0q}K�	��e�����\��N�h�컎��ܳ�*a��˦�+n�0�3�,� ��=Kn�tr!  󆑤-�b+]A�+m��#`/x[�U5=��.��k�ؓ��Ka$@9�˖�Ge�k�ğ�A��t����#���{]�%� �&�[ٹ]+�4�??C_��m���l����g�W�l0�>�oJ�2N#ǽ�1`ó�^�z�X
nx����2�PO�e]�ic�pG@����#ZJ+��<�1�(�ؤ�:��ų�pdH��y����Q��7����!\�n��0�ש��W:0F%�te����2�t�c<K��+a�7م��U���I���8Q����Bkڏ;B�L,�D%M��q0���#Pd�����~x"C�&�?]r�	���ǲw�o�ل��3r�##�h��:����ʇ���2�Å�tȮCh���ԕ�|y�%�=�!ې}��
C���(�Ae����R&�rĵ}���8�M�_Τk��Iie�7bx�����W�J�0�9aLyn�b#�:��Bݜ��2�vwZ������1���DϤ�q?�x�2��m�/��n�inn>���H!�T���ރ�,��3��ȍ����n�laL==�*�[�C___�R;=3#ݢ_4nJ������W~���G{��c�	�۵��Z��v
��I�.��ܪ��Γ<*3��>�{u�J-q���u_%e�O�����:(�=jR5N��[@��.A�KN訃��A~���)if��~�5�jHˁ1rC������ �V^�ޤA��-b�w����]��>�K�r(�1skn0VD��#�����tz�*�GQ�����u�02ͨ5>eI`��4>3�}
C^�G����6����)!�(8�Dz�V���.z���H�Ge� �c�K�{h!6K��Ah�EE]\�"����D�����������&��� T�2b�G�r�7��d�I�ҞTN6��Z)�(+��27�@ ����k��S��.�u�Au�F\/���ߖtpx�vwji{s�4c�7�s��(��D6B�;Cv��}�����AH�&'?#��(�o�8�~�^N�ӡX�BCϘFsĠԆ�.�K��BևQ�V:�{��iS����F5X`��u�?T�[dHBmP��~k�a�ޡ����t��
�y$�z�A	���g ��.��b�獕ׁ��A����,�g�7��	�?8 ~�7�Cz��p��A�x� ���ߴ��j����(�.Z
M����I��j���b�<���2�tSb�T/<ċsDn��F�_����a��N2��/��.��zz��o�Y��-�KIZpK1;L������&��_��v����%B�H���� ��D�jٜ�?o�P[G�������?�����@���3���il��l�0<�G�&�c��)�����-xCgL�P�s�t0�ۉ�9�3��g��� +��R�<�f��^�B�P��>�%�خ�-��Qn�mF��Q϶�03��3�B	F&�W-d#7�
�2��r`�Mt)��J E�N��2Q����q�g��h[ �|[Q������K���.Q�!��2Oe�ؘ/&0��#V�3Ti��r�F(VI��[����rz�Z�}9�n嶧�r~nv"��Ji�l����v��������T��>|� ݽ{G��D�<��e��'J�� :I�t������46�~\}ʘ���+]���E��!fo���J�UϞ��˗�ieu#+�Y�˛O�-)���]�W��L�;Rn=s�z�r�z��є�6>�PWn��Z��Q�-Vn�j'�[�:���P�א�̠���n���h��]��do�\e�ɏa��Ȓ����kx;_��ǄF�m]�)�e	ɧ�c�`]�-�)�;~-��_�׾-ag�a[��*���⑓st� �/#(�0ً�r�J
����Ĭ�I�dF��}o�(moǆ�}f@�� ޤ�Ӡ��O�Z�G ;;�?J�a��^9J�6x�����P�FȐ/���w��Ԙҋo�_�ãs)�'b
�c��m�5���gM巷'�_ �{{��q�)���4�[�r{vVy8$Fe�¾)���H	�M������ ��`�;�/���C��QV������q�d�:�|z�N
CE!�<{{��0�j�xtx,E�N#�U���*&����F� �* �5N��sg�KQRy��8[�g���X>�;��2��S��|��o���VF��N��R�U(��5MJ���I�!{�%(��K��K��,��������Y	@���ܴ���Ud��
3����ʢI�p�NUw|��{a�+C��IRW��H�J�1�ϡBV��X���X�qf�Y�p~����j���d���LSir|,MH��]e�0�kl|<��J(w'�\��YH}C=[q+?�F����ulCv����?�s��6r�ˍF�R:sw����1�ӟfJ���"���~�Ǡ��4B��G�F�Q�Nl���q+^�D�����/� vVj]��S;��SڑO5s�MI#���P�(���!n��JQ+���bEZ���<ǿH?��{1�U@�>ׂ1$�GC4�*+�ƙU��3�/
xQl�}#��H+� �Y�n��g�L�3>.� �����"w�s�9
#J �k��dp��Y؂k)'5Cܗw�[yT�	����&��ܒ
%:�%XA�f�ٮ�
#�<��fVeb�$��J��g�^�t���D}�����tr��~E��j� �Oj�3�~� �ܩN��WF!��ܥ�hB���9��2���@]Q	�!��K��9�����amJƑQ��(������x�\I���VD�:򼯷[��[����ի������FG�ӧ�~�<��&&G��P_ꑮ��J*����Ph'��ϳiaa>��N�q�^&��D[�Z�ՙ����Դ��>)�BsO}�����
���>��,���&�a斛��2	�(���U[aR�AH�5��	�ܞ��r���E(����Q�Xt�VЛD7��u�>�xT(�S\�:�4>fw�al��l�}�{����J��5�9?�p1[ۧE���[��o0hD_��-�[����_��������-���@����P7'< �(r��/�`E1���)3K�ز������^�Z��N����HJL��&�O���\���V��ܓ򧆨�"o;��
bW�p�G�n8=�2S�����=ol��<z�PJ4B��T�靝}���ڵ2ˬ��ށ��p�{mwww�t2R~R�({ �#�P��J���I��%dfca$��r��Oa[��)��-+�ܥ^���W�04�Ueqb;�ӳ봵s�����ҫe+��>�@�?�T*�F��y���"�?�S<�n4
���E�<�@ E_z(W�p �m�o�`$���l����S�ՠ��2LtڤGc��T9U�4B�%�����p�+E�;��</euZ��ؘ�7b0Kڗ�Έ�{�=[+P�8O�y�6�e���H�E%����t"Jr�vh.�=+�t�1�[fmɃ�),��͎I��{	m����c|$�댍{��Ĩp�3���1�3�v���1Ӯ�~��Ճ���:S|ԁꃺ���\�"���Y�@�e�1L�h�n7�h0%B�z�{L�H~y��t�a�P��7B�����E�rA��Kb.�[!�sE���N����zI�0�U)OY�%n�K�9Pҗ����ÉF8�7w��i�K��Zd#r�Xďt��G�g��#��,6`<dcxv�7M��Cy��G�������6�(x��2d�� Ҡa���r8�����8^&�}���ʣ��-�?.*�j�Մ��+�暞6o+���jI��\���!����;����/[q�D���ȭ2{Uf��\PnM��}��+!�!Wf�b딷4��J�g���ۊ���щ-7o�Z]��3[��q��w��ߣAQhd�����`�!3S8��AXyh\���#Ȧ�Q&��]|��	;|i�Af�Y���b;#�:==�z�Q��r���k��L ��?�(�/̤���ԭz����e���s@�a�s.&܉�q�aH2���W�+���(a�Y��b%v��<{�$�f�y3s��"5����j��%�V��Vn�\L��~�>-3��	P�]�6��J�e���J��Sn3�)m�-4��h^��B��S�� GC�{��0�$�v�y�`�uc�OF��-�c=>CDز-�ʭ��r���Wʭ�U�5Up��K���00�SR�Pl���8��5ǵW��;ʾV����O?��4���O��h{{��ﭙ�o�_��"e�4�x��m)���4т�a\P"ܘ��x%���2�%{����q��g��߲�c=����Q 3����n(�uۄ�����*�'_!a�mM#4��c�P}��
��P^,xس)w�������F�)���_���Z�X��FZ][I���j l-`S����3+���ח�\F�lG`����\�ͭ�����^�\�u%42fs�'H#�[���%`<T���t��G	�������d�a�F�#��r�����I�c0255n�4;7���c�/J���6���,A�):���Y��x���E�������胻��)��R��?�:�V�n~z�Q�k�����bӕ�l���>S[9:Ԡ�:���ʥ��N>��3>>��gz��������3�쿞H3R���{-E~PA��6��6��!��7ƞ�a�Rp�](�lM`{
{����`�X��&�n<�@�d�����`E�,�S�7���v1�3�`��MC8|��Ƒ�54c�9!;E��~;͟59ra"���~���
n�y�n�O�x�
�H�HG�����w�ZڢgW�?n�
h�'���2X�A�u)�#���@%Qm�i;�)��/�S�~Ȉ
��g�g�r�_��{����lWϤ�ethPn1V�=0���t������-l\�@�x�uS�T�巌�Y[V�P4h_���f= ���~��)�6�|G�Z�CvM8�<!�P�P"���r�BN�1�g`+U�,���4^R~P�8�6�a����8�<>���]x�%O���	{Bx��Q��@}�x�>��5RB��ݴ��x֐��/~��,�<�/ ��]k�P��_L����¼�#� L���Aч	6&HPjٚ����n�wo՗�ׯ^�o�U_~.:��{�祐]50�D�G��V?�'�|�k �/�ؖ084��G��aZ�_���YѴr;8�&���G�)ߦ���r�:��n�r{q�CP�:�[���B����A�[��3���?�'��ek\ٖ B�s(�����wc��NuQ�+h��L�$�n��Y#��r7O��(w�������9~����?�f��z���6+�q��]�3'D�r�����[�$l���}ϭ<c��y��3�#Ǝ�ˊ-�,��s�L��[i`� ��'�\0ՏO~JO�)=�驯�8�0���Nw��q�dF���$�xQWn��-�)&4�H06L�V�8��B���d!(v��?��<-/�x��%}�+��\�`6�P�>��/e_�칔ʸ�������i\���

�DF�(��v�g}m�`_Da�/a��I��W�^i�k'�����b�:JN��i��眀3S����ʧם���e�ب������k��+m�-�?�V������Fq	p��CfǛ�%C� ���
U��f�z�\Rl�,�/hČ�9?˵m�Rp��qLM�a��2:�:bluڜbeC�ںd?���ˍ_u/tY�푐K��D�Ό��;ŗ\Յ ̸��L4����}+_-��ʢ�൳�3����N�\_O5	�IBeV�Jib�ݢ�؊W�_���ַV�'U�;�3�k\<:�m
���.��loMj���]m>L��w2�3�.t{��CB�K���p�Hkk[i{k/J��r��2{(W(E�m����wW3.3e��)\�Q7z/������)�p�*B@�Әn�x˔7"��-&�;���+��H��K�Y�N���$h?Z6'�<�]|� :�*��)mQ�U�2�[$��
�N |�o܊r([�nsD��YP�o���6���ِ��^���<�9��~�9C1ƼD�4�4����p&���ϱ�ˊ�A~fN�ѐ�[�<��.k��!P�SN#�5\��2�l�c��uhx������Lf�Ќ�+��=�Bˍ:z·��J�B냿RjQp��`MJ��4�rs@�{O9�O=�~Բ9�~@Vq��4����cأ?=={J�u�|8O @�pa��3��4�8D0�]��]��+��>�*,��c�ط+ � �+�	WlO0���$�zD�����S�%?��P^�_<�K>\�y�z�Ǹ�RnQp�( }VG�<����j�g�b�U����I#�������![�$b��LL����������ޭ�ziY����42� Gʭ�n�Rh���iemӫ��ͨ��m�Y�{{u�z�/���G��Rn���ʨ?�	�߰M��<1e�%���gn�g]�2V�!o��<���𬴗v��!�9���~�w6��_�6�r
���6��y�,cUVh̝�(P��g��ܖ{n�mHz��5��D�A����������=��؎ ��0F�̌Hȝ
�ը¸ѱ���겦̯�l���;�����9��-���ӟ����ʫ���� �H�~��Gb�i/��/��󵴾����R8���	�x� iL��2c̒��w���t�O~|�VW��I�f|�wI8_ECK��D�d!��e�|r��D5�r{qq�<QXQ�84�2��FZ���ݯѵ�q�o_��""�	��CA��yv;F�R��	rsa�=�R�%|F���	�7�&f�J�ъ+L�K[�r��~��_o���^z���'Nw�� �q�A5�2�"�궻��� 3g q#�.^��0�d����]��lR�ǆ<¶�G����s�ff!��q�W�AK�G㚖n�e��NR�I�?��ȃF�^ۦt��O�ή�44�-3l��V��Ĳ=�c�C]�3�j�\��U/�H����A�&O�n�I��lX�==9��> �P�5�kf���$����Rid�F��pHVn)״:D�D�ѓV�Z���?��[�sO0��~<�Z:	��۩����Rh_�^�3�޲��)zڱrK�Ȯ�UU\+�n��k�U�?AH�� ���_�{�����T���S(�b�V����=#Pvsz�WV�h��Jt�Q�"�f�?ʣq�ԁ*��v����p(�0���u��A}����CP�YiK�_)��)l�e<�!��S)e�ޱ�Tpl��[6���̐��]78��?l�pr]��"ٕ���|o�mA2Ge�>��Pn�{Ňޤb>'�W���zG�ٿj�AKِ�n�圄���\��J~ЇMό�:�?|�x���d.��#j���hzZJ��1�{�9���~yfkǥ�N�rE8�A��K�k��l��C׻�.Ifp(%��m�����\({lOݿ�t�y��ޝ9�q����ǖ��������/��L/ڞX��Fs�3�'��_�jO�|fV2�-W��ƞUG���6�X�Dn�d(�AQl���"ġ`�0�y�%��?x`�A���#*��*�?�E�d{(n	�$�0*%Q�mKsR�z�'�n����j��ܖ¹/�y�:����T�ã�X���竭�O��*WJg�A��e��;iM���ʆt�)�+��K���'�|�T���>L/^�*��r{�HO6�n��ib�C�33Sq��A�d����K\�M+�b��q@��<��K�[lcdU�Ʋɴ�6@8Z+�z�Ng��w}b�7�R?�e�m�6s�zop��J)�BD��$n�J��Ed��۞n�R�/r�ʭl�(k�
�w-�����vk;�ۣ�!�,���Tn���tAC(ـ���`**�)��;w�5��F�>F���{�P��v���FQ��) wӧ�~,��P�io���?�v|���(�e?p8�h�@�eK@��e?���G�ɣ��O_���mU����z����QB\�o������p
�=�̜�}�'�E`����]1̑�+%�S#-_�5�����1_f���{%��	�7�?����yf���Έ����>b�z{D�)19���*o		�)�����~¦whx\�T=���͘�=>��{�c�A]8@1@��&��_�~��@cw2r����	�&yK�p�X����=����}	�������/� ���1�L�ƹ8�o����I�\-w�aI��hN�#ݞU�^a����O���߳��_��������e_��������K�l念o���%>������A��Z���6�}�oU�M��NZ���]����3����q�"'���r�f�#�L�s����	�A8��N�ig���!!_���F�=(WµY�%J-�F��y�S)�,'�z�����m0����gL�w���8��W��b�gY���c䯘�W���ֻߊ��1a"�@'3�	Q����  �J�A�;0n�BiD�tg.>Bv1<�>[���A�H׊��+��+nr��T�Djo�Ht�p�a�L�x���,/��m����%�g��o�3�3�		�·^~A��$B��r~N��ɧt��q�%ۂ�Ϩ�$���.�!���J�]�3�~l^
Ҹ�{\�LgU.I����[�t�~��~)}�7b�;��n�vO]H��l���-OTx���Y��ag�V�[�<�2�@|���k������-�4�D�JK���� �/>g YH?e�3�7l�_���|���p7g��gIX=b5�l��\�l���z��E)��;�G�Ph_�X�(n����R��*�^�g�ߙ��u�q3�hAݳ�o��
)���[�X2��|bŖ-�{i]����
c��R���?dK�kJg�6�'���^[w�瀙��h�C|q�6m�I�]Q���م������Ly�3�L�������";Tܠ��١6C���zcv�3���j�6>�A3����A����ꖖe��M�s̦����6��춬���ݣ�	�#-� �nu�z�����_���S�eY��+"[���m	(��;����_�gVn74
9�H��9(
VnK!2Rk�.���LO�0��TŰo��|әwf�@_}�g�jM0R�V����4��=��?y����es��<�2��6�w5�઒�;���Q��B�,,�H�t��ClK�*����咕��N�q���x$����C���20��=L�C�n�\����*�����ZI�M��:-���<C+���`��J[e�.\�477#�uhd�E��΍��(�A_�֢���#)Z�R [ӌ�[*����p�ܪ�U^�ZV�S7��/����2kR�q�F�e~�{H���s��?.���gVn��`�H;�ET/>LE����%p�*���)m �fqp"{��4:�\H�"QN�z�qs���c5޳K�?f�ػ}uͦ����4x}�T�=���%���Ԉ2~R���Ex��nnl*̚
�Z+z^?nxo����FM����t4��h���ْ����M��.>G��J-3���x��)2`9>:H�[��(���JyF���0�A��U�Þ��MwB(���@Y:S�$|�n)���J�eP(~��K�AYRg1#���Rʭ��;�bxnx��oA��Mo4��'ѥ�����o��1���7#���Ļ2��JRE��B�Ep��qYr /�*!k�ŖA27�"����L�['c�aď=��s�[�KQp��l�~����]���3p���E&�n��T�J�w���M~vG��Z���P��l��b�[Vrst����I>�γ_�5v'L�s���bG�3��r�I��^)GS#R0ƤDNx��&��M����c� �-��j��~]�)�E�\������$ch�g��m��+X�b���Ӑ���,I��-�XD�e�=�+Jd|0B �Ϲ����ɢbK�(�b��$Z,w�v-�ҩ�CFB}#��������D��<��l��t���~c���<Y�c�Y+/����Z)o�[�q0�7��a�����������X!�`V��{[���?!��^/��5��r��>�� m�>�֥�.-��G޳=Q���(t$�R`_�x���R��(��Q���'|~��x�h2s���r+�z�m	f�q��O2s�~���L�p�-{n9`3��G�U�ȡ+)�Lı��J��"�2�����:��oK@�姸n�2Ќ�I^���R�9���;Nxb[�Ц�A���-፸��i)��`]~Q��A�u0����JS>d*e/�����-p�OC��C���rbΜ|{�Sܪ����&6�r���̼���U�61�YO�p�l
ǔ�G�_|�~��ߤO?�,ݽ�@#�~�r��O|_���s�g*��X���j<��v4X�Ro!\�h�`�Ң��Gn��h�R��`t�e���^��r�o�a�@+�|�'���J�0�G�i���w�z���`�G�(_�%ŏ�o}�5JK�L��L�en�ŝ�8Ħ����FK�T
G�Ja]�����h2SU�;��6
��A���24�޲��\�3A�a�5��:5=��~��E��O���_?I��]��wߥ�����_�/��6=y�T�����؄��\�-!�)��IY>�Z@a�]:W𢱠�!���g{B�ẝv)�|8��fw�$�!�!>��Ԟ�U���fu*=������4;5 L3S�iz�/M��f�K3�\�=��gG��4_�HC�]�L4_�99>Ԁe;m�I�-K�^^�p]�rʗl�D��Q�.f�bi鵔ؗ�v
Fq�� '�~x���2��[�Cƣ�Ͻ߆?`��y�}Ƽ
��\�P�n ���!c��p7�W�\r�[`�ϊ��=��iw�E�?3�f���ԅb�r���o��%�<�/$ ��?��N����W��}�(���t��q���JP�;O��dS�7j�!��R.�D�>ޫ��[A����C�U�x��W-�#�W�Y�y	V��=�4������������Z��Xf���A�m>�7�Ӧ�m�������P�S����k�'�� X�Wgǵ�K�7]H&�����V��_:S�����$Վ���zZ_Y��x-\�ZU^�Y��&��4[ �����!ׅ���l���j�̔W��vV�$��*��g%��>~x'}����٧�ү?�_��������Ƀ���tWJ0,�W��
iru'^����������ݽ��5Cۊ�e�R}bJ�hW�G}�rS{䳹���KKRV_�g�_�g/��,x�,l�ٗ���(��]Z�U�̐�	^z!�E8�@��f~S(C��g��Ɍ� �s��]Li;Ya�?�R��J(����u>��h0r��'@#�s��+�<�� p��|H�1��&g���r�r��k��Ɓ|ޤ��/�߿��=T�:to;@�8t.?��Hy��H�[<�`�z�ʑ�a���׳(%nD��I���U����.���LC��U�Ѩo1��OJK��(�"��l��/��+��6�-12F���t�\Pi�C�F�ܺ��Ni����=5�a�䫗�}�{����Ø�EUc���	��g`�{DQ�:��R�W�8@���sᵣ6y"O�  ��IDAT)�./C���=�(ǌ���c��=��8<���;;;Q\��z�%F�\ړ`D�p5$[!�9FѦ�/υ�)׃+��ؓ#�؇|zz��g��.-��jNm
f�D,/i��Y�f�p�A	?��>�=\���
�
�lo�q-{��e*}�ɣ�=~lA�pַ������7�w�e��o�O?=KO�><I+�˞���s��O�8fn�4�aՁ[5ز��B��L�\y���!� @�73��\s���^���B>�<44��c0��i���F�|4�AA�Rޫ��W]���qc��;���u���.�1Kۥ���R&�>��Y[Ǎ�A���t y\I(��7�#��@uկ�"W����i���v���T��O����m	��C������o�����N���n��!F�BT%���&��W�w��M����Ǎ8(l󐟔o |n�>+�h�?�D�������J���ڪ�J�K�B�׳MVD%k�	D#��$���L���N�@tBzfkc���B ��0$wb�6���U+]�`�7�܃t�)�_/�0%Bq����/�+�f���@�xϞ��K�"�W�YcY�2��;c[:=ی;�\f�+���_d����,�����w�Sv0ҥ�K�\�>�k�q�!��/�s��x�"�~�J�p%V���%�co>m�>���oX�67B�Dݔ���o��߸�]b@���c-�܅��wd@���8��
%���>��t��O��}K��){Symx%��TGG��N�7$/X��
�����qH�/n�L�\Y�e{��j"�O?Ȫ��?�����Ϗ�i�'����X��J0x��������!�Q�TK����3�� ��$��[R0��\/*k<�x�ٶ��>��`y���O}M9L��-��㹾�e�d�C
��{�K��+�{������/c+ة������ܢ�
 �lq���hS݌������4=;�[�]\�U<����u!�=�$7��"�o�T�-^����J�X�A*>,��j;nCj7&�̭�����S���Ev��tfv9�t��l����`r�L��4'L�iMK+�A)�4*��l�渤m�μ#'�Τ7%PO�ݙ�>���~�-AeFW��ê��`��R�u���gL��c����&�K�D�����ɫ���Oҗ��>}��O���%5�=)4�!=,�B
Kߠt�v5�c+�?=y�^>_�R��,K?��d�I���,0�"4�R�	/0CK��C���tȍ�Y����L�*�5eFT�O��d�;��ul�CgŵP0�i�����R�2_�Q2"qz��BYGcD��,,�������4G�fJ/[x�b
Cљ�@@��2U��ټ$~l����#�J�1ރ�UU���E?)���]ݖ�RNϼ�����!}�����g���j��,�����LQ�}a���	{#6�)u\�����>ʰ�W�GЌ�Yާ#�@Ug���M�K�=����7�qBV��K��_�jLJ���h�b:>:��&����h�����I�c�ij��Z>A=d�yJ�~|��t{|{<��r��?�̾�~������5�oG�_�a��}�܏��\^F����Av�~�����ẋ��=�x�揽�#M��N2���b�=3KU�������Mɻ W��u(n��iNȑ��zKm��@�8�2s�N�t*9�b�8�h��/p�$ekE[u�9u�V�e�=�.P# V�~�	LnR��۟hJ$�[�N�]U��$�=���ճT�+�a�/��q�� r�(����1;��[�T�(\�RV�h�<��ϲ���Jz�2ؖ��a�V>� yBu�����mI��ܐr��&�v5ՎvՏ����>�9s�R�P
{��h�dC�� �z$czӴG �qX�]�VJ���~�C��X��3�l�ڗK?R��
8��-��pK�>��K|���aﱿ���U��OQ��������J�����Z�]��!L��[��6���{w���;s*3T��"�3k_}c?�F�#�QAnc��^��@XC�}��X��uY{$K����CεLLL��6�s��C����]*u�֓��3)�꧕�z�{����U����P��$�=�%9�hBV�S��9l~�����?r/�x�w�y�������-�˯��� D��~EK�ѳ���]� �/���� �����g2t������
���+2�H�T��H �3�9C����3v$F�'j��v�?<I�������W����������u�����o���W_~+��F0q�#N2��䇧雯�+̓R�ے�x��'����"O[?S���Y���J�ef�����bXF�*��Cŷ�����o���ˌ�g<J�r�0\�\�`BC�~���$,؃��Ŧ|)�5s0�Y*ß�u�G}�)�#%fy�Ńb��:7َ#�.�\�`�I���T>�R�`��%�C��2s��z�3�@�h�fb�:�[`�&XYl�@�懝��������WRH1�3�m(R:�$��Rf���6�Ll'���ɩF֗1���F��+IH���j�֯�Yک��Z�-�DOР�`��Uf9^)m�Ͻ8e9�ڃ[LM�KI���0����^0C��˶�6/�wHq�2�#��[�tڿ���˜�P<� ���4�C�YdZq���2cO�+��9�`�1��XoU&��hō	�= �x��m�N;�䆩�i��!��^�K���B��z�leS�c<g(��8�*�ϽW��S���8	��ET�m��m	�*�PnU(��)�mNmϳ��{+�����2 2�.ĳ���ˀ�cL�r��!E҂f@A�*D��iS7%Ne�K�����%�k�!�3x�\��:A.�+��=~��|-��{"��0k�F�+6L6�r�D�Վ�;���Gi}}S��g�Z��(�q-���Y~�RwG��7�V(�LOU�����}����G����Ox7ݿ;%eq4-.�������x����Y)���I��<��3|�wwƇ��ߝW���gK鋸���ܳ��ˆ�i���"����m���!YVѳ !��GY	P�)<�d��ۛ�$��^�����}|qc�����w��}���O���!}�������g���1��=�-����r�<J-���E)�*�^97��/a�-�(�L�� -�:��j��<97C�9�8�>��q��g��_������*��ן����駟�?���-zv2MN�{���T�{�Nz��������?��a>|����)��57�f<Q�`D���\�����A�ɥտ�D�x$��:/����r䑡䉝��� <��BR�Z�L�^6��|g�C\�<����@�1�U\��ϱMq?��igA��XA�A �9p1HI������|�ՋW��OOӏ?������������3����Ӈ�Rr��W.�yS�f��g�(;�.�#l�HE�w��P7���]I�Ɲ�jĹ,�"q�(��%�X�/��$׬p(L��),)�J��~\>���<�0����{B���s	w���̐z2���������AȳGBfdtT��!)�J�Z�31m�"Aӭ����zopx���Rb��'���eO`��7��&xK~j$1�e��TX�,p��o@�{�a���)w�W��̏�����?8,|�rݕavЀ���@��,�p��\o�=
MDT��1�j��|����^f�
z}�x�SЃ>����%��B�r�(DG{S+�CiR��.l��A��NA��׾�H��B�8�̌|�� ��ɭh�����)���3��b�ЀG�ř��av������
W��IA>FZ��KCC4���(_n� ˣF���o9-+m$�@!�bW�+�P���>�a�^�9M�G��W@�|�-�N�C����P�����'>��eP�4�iw��(�Pbr����H�41ة�)0&,J>JB�*!��i~ƁG�1��p%�LP�$0�\��(�V����Q�u�
O��V7��g�������S���+�( Qrx�*����.ŉ
2�<�=W��H��'�v����l�=�fq�VRU�:4�涛ab���icM�;�	)��ދ?39$e�}����)����tHIm���!2fBǥs�W�D��|�թAp�p�	Jig{{��Q���'#�&��7ԅI�07Bg"(���?���r�ʪ�9�ig��7}������?I_~���>7��W?�'O^h ��:��l��|������-ߔg`�+u�:+m��}g%�V�Q_�O=�U����I{��Rn�.��>� }��_H�E��e�կ~a��O�g��8��Jq}�=��<�+��>����������V�?���Rr�K���g���{r��3���v~�yg��`�f2�>*C����ʊG��-���^�P�#!�9� Ф��6(p��+m�.�2'� ����Ew�w�����u���O%��1���Ա�+�6��g����~����`�,�'\c��K����g�hj�wl�Em�?���Vs�a9��yf.����nZ��HϞ=O���������_��_�����MO~�!-�ė�8���
����I8�i����y��g0��Mq��]Xs�rU�iQ:F��1�d�Y�V�A�Bid��J!�)�g�.C����\�+S�_�S��H`���O�vtJMC��HI�6f�O5Re��q��0hK[V���Uys�.��eb��M����?0�t�流1 O��zc�O���mfPY+л�c"ѹ����4���)�u%mR��%�h�� �=s����^��Ճ����.Eׁ��t�����Gi���469m%�OɎO�h��PB�W*H�P����j3�|�&�:�^�v)��=]J�:Sg"�ɒR�p�����}=�	M�^�	f)2��k���(q�뾸����%������;T~x%4�� 8�[��\(��]ɩg�b+oI��hoM)��7�[�#��ON�S턓�\�,,ʌ�X ��.��"RU(㹝T[����U�4���y��ޝ=����n8��07��H����!-Q�~�8�D�5:(��!eS>W�����	�)�12��P�;��L1sX�ZP��(�)�j���=eSg�8�A�Ά+|�;9�^�ލ/�6�B���BF��2e��;��)]�}X2�*��-��)� c'���#e�̀���dŶ��?�q�*
ڸ�[���q�r&��h�&��#\
�C����<jw(U�
o"�Νc�#m����{�qGw��N�w���3�Α��(�)�	
F����x���Y�Q{}�&�J�O�M�.ĕJj#�_�R?p}��ܛ�FF��L�A;99�������S��=6��z� wۍmN�C�^	��iN�]M�[�ߙ���4=���we�U`~vZ��7�H�uH6����fjdhHʲ���!��U&)-���Gn�D�f��Z4�P�=�"��h�������՗?���|����J_|!��w�J��&}��w����� �*P}k��>"�|�*�(hW�<(�z�.�/m�����&���'E��o��e��.�R��?2>���[H�|�A���IA��'�W��XJ*�I�3)���|f��?���_)�����a���/~e���7�/��/�?�'i��g��>�<cN�R�� +����ҩ~�iS)���
ס����G�[Uq�H6��r��3�j7�=�.��6�/޿r߁���}4�҃Ihg �A;���g������Ri��1�X�[�B�09=��vd�M;4rԝ�U��.�,Oe㭠a�r ?�c!ȑX�"��6�O�#�N�Θ@'���p�4��3T�.e��;]94�����\��4�����n����iM
^6�#����_o�C_��J�@��M��,�~�.q�+�(Et8�lD� �L��D�EE�0���]X9���~E�K���:�ސBR���-��T�����3�\q��I}++BN��btDE*5 =���P�8Nɋ�:�R� !�F8��Y1.SUnޱ�b!1�g5eǌk�h�lLpl��(a ��#3Dz^~�%F��1fI���,m��H���!?:�{ll<�W�����_G��H�S|��+�ަ�����ZZ^�H\�EG	j�/�f�� �"�q�ni�@!����NgȽ�q������ُݮt}�5y�9�������	<d?5�&������D���3��5w�šD��l!gp�\�����@9�G��W���lc��);�6�� �+o���|�_�$�g#~�o�JXp��3�������q^�s�?+�%Zv���]�H��o����X���	���ф�v@�gƦ����e�<�ʘ����F�'Ӆ�E9��&^���-ҋt����˕���\�r�W�G��'G����ov.�mJ��/�)���򓑓Th�-@�z3OEB���b±���P����F8f��ʌ9�Ѡ;8S�����^
Fܹ���b��\oo���a���=� �q[)2ܛ�4�J}$e�{e�ۓ���vW��3�-��S
q�o�aՎ���9o����*VJ�7�0���T���.�G���h��D�P�-Ϟ�)���"e�E��6!�" y)� �B)C��?c��@J���~Z_���ݴ��#�J+����ʗO��=9��D{{�ҀO�N(�y05��P�"k7���j`m"�;�T���09�P��>��������A-�3��<O3f�� �����\ [�Y��?�0��ĕh|6����5}��7����#�ѧ�@D�s��ʴ���Q�e���v�|0�O�V��C��P;�3�·��a�'�����=�-7h�@���<����n'N�!� ���'�<�&N��<#�,K����H��2"�?�4NLo#v��/��N<�n���N�O�=xp7}����_~�>��g�_�>���������\���L30��aQ���{�v�#�Ï>L|�AZ��\���ϊba�՘(�ćߣ��NQv]�t*<��� bj+�(�w:��b,��F(�R��
	[����3��j(��흞]���7L��=�4R���ڻ�^�ph�B�{}O.Ҿ����ۉ���{y�ˡax�1��_+�����p�;@'�����|̊���ИU|��a��y
"���8anG�����s*��4�+~vR1C����g�Ql�bp�z��p	6�vӹh�{%��U��h%��{T_�{�|%�z��=o��f�%6_�HVf��g�d��l�U�1���M'�I>�p<��!Z������[+�\fw�*���s�������D��L>(��ܶǈW�IX�@!G�3�fP�a1�w	�J�)}!C�CQ��\�+ l<T�@��w�c�;��S �
�0��ۦԃ���P%��w�y�W`�i��"�e�@'xWy�]��?hn!��e,���eep�.����6xSc��N�e��ֳ�����Pr%=:��g��tLNKv}��	�$l����s6�7�*%h�m:��3��Lkp6����;�sJ�|��p��  9�_bc�F��o�ߌlΗ:��B�Q�B8|#����
����/��3e�DL�jlK}=ܒ��*@�i�q�`|X�:�}�r˶�N��qϹ?�-9�do��)��~��~�U�����~3��r��+)@d�6)���V���NO8`s�$w�����1p���C�ƶfh[ؐ1P)��\a[��8� 9r<�[�Ju��֩�N�k���ާ>Ԧ ���'jk-�V��peP�~׊(q�g0d���T��8��h�ñ"�&.j��R��i��=Q{�>�
�Y@�B�P���F��Orߤ�kP��r����C��6N�ZEV�Ӥ~�J��q��;
W8ѯS.���Z����J���~z����C]髃��n�5(|���������{D�����p�&�g�_�~�|��˚1!�Ɩ�п���`5��K���v�
6�$��A:��P7���� 7qȉQͽ��Rf�O>}�~�돥�~�~��O�ǟ~�>����|�ɇ��_H���a��p!ݻ7+�x6ݿ?�o*�O�[������?=�mT=[��/�W� �.�q��U��Ҟ��fcV�r�`|��m:�ҹp�vPpe3�:�J*����v������u+.ڧA��Fu������A�ΡfnQ�4.
�ON���HqVzgg,���ʭF
^�C]Ql�'
1�K���B]*��na�i�����	�c��@�E3n~���2#��r}!t��W���ZN�n�oV'vOO��ۙ��@ǅ"^J�аH���k�58X[�0�'�B��j�J��X����9}-B��cEI��H(�~��j4*t%,F�UH�A#���@��)hy�t����G�r\c)>��)S��Z��s#(\�e+�a��n��4d.�����D$|��UH:��1�@'��IM��TJ"�T"¯3���[@1Ĉ_���o�9�H;:���[����ߡ���i9)£�Q��������@ϱ��((���P����	�'�S:��E9�@ݟd.�\v�4��}O�+X��V��@�[=˔�u�H��&�)��9he?p'%���p���v�z��%Nc��D�;8���/8�l@����L��qo/�)���A'�xՃ�P�(���0jQ~	���Qf�-V���2��BI��;��SW\�%��\��$r���$��;�8䲅��$��e {�v@)��i�Ցq�W^�R��
�{���pY����K;@���3�6g{WX�r��ח�R�|Y&\�04��L�=��������/��UP�HHng�#j�=�XP*��^�CY�	Ź]y4�?��]^�J��6�nc� _f=`�m���{Sa��Ӧ� m����#�V�����Q��!�nl)��Hgu}7�^�N����ʦ�w��Q͓Y��횎���L2�������J�(8����E��ǜ��4 ���i�&����\8�풧=�'�f�/:*pү��ȉ����{.� ���(Y��k�s�o#��v�u�X���llGfaI������ 3Z\�126���Fӝ�S�Oӧ�z�~�矦���ߤ����O��!�/����y���7�_����=�Hw������9�8U�h�������[�k��tƓ�{�,���Y~vi$l�6G�L-�x6�[��m^�C)��b�+�����X��D�:�f)�j<Giy�Ƴ�VVw|���2�B�������rs��7�T��S�Ԓ�<3�;8:��ˬoS3�x��1��А`7I�~;>�JA`�P�bY3���N���c3T��0���G����#���}@��	�Ņ���0�gf#Ԁ$$|�jZ_[�59GG;�mMAO|O��w""�v��|�p��c[�h�&ы���%(Ԫ��C,�QÌ�Ė��}h�($ ���	��e���y�o�l� ������_eFh�Q{2���
T^�Q^�a�$�����PV�;TB
������(K��? .�_@$�c��O�[��[6������e���2
�������m^�� zˎQ�����!wvY�j�<|Y��3q�%����,x��+D���4�����L�?�A2r��].�E�E1�;�B���.�GV��D�����ܱe�(/J�ڒ��nK���i�(c(�q��+6�y�S ����q�%�_��3�D��rȲ��cz��Wʭ+��@g�b�S�4B��6�/��)�ؾ�g8ԓ
ȿ��y�zE�m�J�g��5{�ܮϼE�é�3f��B���n�1���qXͲ�<��~���m#��A1N�{P.��� ��c2�{��L<����.�}�W�tw�l.PT�)���0��Jf^�mR���R�v�j��֑��F���D�J0nk��0������461櫲�r)��׼M�s+Э���y�(��B�ۼ�>SB�S��i���-�Kem�.W�\���U���g��_���~����U��K�e��W���?��E���_����_�H��<�^�~�����w/��߿J�� ��u�����շK��o^�/���_*�����R�/���I�滟ғ�^H�]�D�9��"�8�:I��L;���E�4#K9��M�Fw����(��-�v�Az�Y0G�Dt�h�����ŸU���.�[�SUri��/� #����`g��Qz9M�s\�W�@CXA���mB��s3@d�b�5Z]Vp��S4ԗG� 8�8�e��[���=93c|DṠ�l����,u��rG�U���XB$�9w����<SPoL��<[�Q�7��J	���Τ��O��w��b�VJ'�-�h[G�q���	����+���i����Q�Fp<3[��zt,�|�{,�L���1��Wi����L0{��v��� �F)ٟ��#)�R���Ga�}+h.�L�&Cf1��XQ��i4&@�^�$�B+Ló�f�!��Ϡ?�%�Lo(����G�f�e��1�ײ�:�̫T�|��=k�4����|��������|~W��'Δb鑡 X��(�A(��6C�cV&ff$\�x����)4��\t<lIa+
�;pٹx��-f�Y^R�Nd�R�*���-�k����U�
{������?�XS��4�9���>H)�MocF}��Z���þ���S�����4rZv
�*��A���{��u�2#�{�%z�~3��"���mS=\�f��ɌI�0ؙ�7M�7����4�!\��v��LpW����x.�UV�+!�*|c�6�Z+��I*n�+�9ٸ�a,�9tz�g�,�DZ��=��CIC@�ނ&7奐�&���K��)g�h����א��6a�8��ܔ�өL������3�^�K��6 �D�8r|��� ~�\�J�ң�n2���D��bK=:O���|_O�j ����Ftd�i��U�(_��D{B�p��e��Z�iȨP��ڄb��7�x2ԳS����pw

��,E���S�kL��5��W'ꢸ}�ü��](��	��z���Ttnb����?lqxx(\ZiFy�U����he❁2��[Z8x�!Z��O>�ׯ���o_���z&�6��F�R޿�2�����w���Rj�������_�oxi����򓲌�+�˯~�R�D𣟿������<K�^��gw�:&u�t��r�V�I~�5�U.o�R@S?�q��J�ޣ�U�*����[�Ÿ�s�+m��.Ҥ��JM�p�׍�T��'=�U�y�cr�%.ab�8�:��z�^Hܑȧ�+`w�1D_Eo�0%`�K6�p(�����f��srz�VJ�u::=O5u�gR�.�����բ9��(��H�½˴�s�vd��@e� �F�]铕�#;�8�=F��ad�N��B�#;fHB  ,q/(�A��n��)�x�İ�e=�m���N�C㩻wP�v)�[)�\v������s`NJ���sB��=����q6��O�w���4 ��m(�����>᠕�?�L�R�W�v����#/�W{wD/�#4'�X�E��=I��Ƅ�r8r�t(�{/�������˳�t����BPP:zF�B���v)�#���铏?I}�a�w�n��O��\�=&�̤�Ǐ��w����TZ��ݻ��Ν;iva^���?_#�����;��PDC��2����f/}"U���(_"CyD�!��g(����bv��P֬���|���(��CF�E�mM�Mm�v=���Ƈ�/�L�O��{�~���w=s�Á�Qx,yr3__2J���n���m���s)B�U
p�S�Fw�S��r�O�����L�l��Е���0&�%� �Q~�#�G�_~��e�{�P�,LB`a�8N����p(��`��0�� ��ӭ��V���6����rV\P�B��^a7���M�;�
:[� _�D�W��l�&y���u��a��़����.@�i�9� �v�/3���'+D���}2ݝ�gY�3�q�J�xw��e���u�ʘ�@�?nJZ��D� ��r��U�j��)�K�?��:������/%�H�RV`ꦞ[QbFK��'���3�KڈdBBF0���`E�d��Yr��1��v�Ke2i�
I�Q�cebZ	�X�#�"ʙ"R]��Ye)\��¢|��YYJϞ?OO��L��V�����S��p�C��[��0
,���b�O^�~�CN��m&����hZ^�5�D?(�2�F��S�)Z5s�B�Kh���o�ѡ�������j����Rn��c���'�)��oPH�}*��i���g
�"}�x?π�3������7�F�o�Q_K���+о�b���'�G���땴��#ٮ�Q�.��L��p��<��bRoq�3�����P��n[~��28\��5�*�h������T2� I(�h��?Ř�K����n�)�X�6��.���M"Ռ{���?�Yީ7�)�F��p�X@��Y �S���"s��`Q���٫y��륭���Zz�rE��`��/_eP����Ŋ��������]}	�j�;���	8���F?�6~{�\�/��iMr��ƮF�{is��J�{TZ#�J��!��%dw��
+JLk{wjk��j�jHRpρ� K��z�@b6�Yte�m1닍�L���+8��Λ��mln���u�iU�d)���s�|�q3q96
�Jf�xP�;�Jx7ت��n���P
��!)>�ө�����`?�p|O@u�O^|&�J�&�2#?>6�ff�|�����lz��N�����>N�PJ�O�������4>1�&&����X���wU���g��g�<k+\�i�y�qƉ_)���L"��ʔF�����OK�=<>��:��(�����k��I��\(�������,��Ǯ�]�{(��W�P��wx{�T���>Q�"�t��;uv�}���Pp�c,[#B0��*�Ȧȅ"H0n�1�L<{�܄��UA�sۃ����������!�r�ü�PGY����%���.�@n.���)���X��k����o���d��dP"�i*?�1��0�����ue"���v�c�ۥm�e�u�Sʻ̪*J��P�
�2ƭ!��A��R>A��ˋ�t~�^�W�]�ʘ(��E������������qW���R��6�R�׈(l�Y�o���Fg�Ӳ[IO�\oQ��n�D�E�S}�G4�B#fE�{Z;a��V��^b����ck�+.�L��2?�@��C��'�E��b�v�A�A}6n(�я�h���W@�d�Y6���l.u��(Kԍ�'Ӄ�y��;�v.x���ں�u�SےY��P�J~V�В����^�?_^^��667�	&W��Y��l@���6��U�
 �g�> P߫&�!m��p�k���k;>�������6�q���o��^����������np;�acK�[�[ے�{���x��z�8�(��Z~�E����� �����\��
�����{6�1B�!m�29^�Q��W耍a���3�=�v$~��ݖH���HV�Y?1��\�!?��x�[A69��n���4��D�xVD���1�E��Na�Hĉ�N�1��QH��HI�򷲶�~�����/���÷�o����w�����ߥ���H�o~��ǿ���7�w�{��B#�o��>�'Y�(���,�P'�PPJL�����@a����L�I�)�Ǩ�����O�i����FZ/_��һ#���_g����⚓�@WT�1+_�����+��kk[����B�1�l�"{*���]i���fZ^aO�f���(/����+�����u������o��߉�����wjD�R�kJ�ZA�G_B�!�$��4+n؂"�݁�M4xo�������Y�N uW�)�݉���#����sf;��L
�<E����w�;����;��Ï�?��O�_��Oe�>�����Ἷ����ۛSo/׃u�Z9.G8�,4��m(��M�%B�3�I��3��0���G�p�,u����~�g�&g�R:��N����	�}�d��Ҏ`�%U������w�6w�3;<�Jq=M;�i�0GJ��2��
O���yP�{�9�x)�1��ٓ��9T�)�ڄ�M*���3��/��\@4Q��u
[���*Znն�/���s���5@1�b��AD�> Vnŧ(?�9�8��l�%,T���/�C�m+�x�#{�Cᅂe�G9ŏ�$<���&QBPVr�t+f���J;��ƾg�r|ˈn.h؝A�K���E��c���s��r#�Q�U�	k�Pʐ�[�Wy��|+%Ġ<�����4������Ur;�߆�_�D�~��6aZC7�ū_���OР�����P!f��(��!��R�s>���|�
:�أM6����/��=�]�pr҂.��y�W�E��q�4�989}\�t	O��m����^|+��[b>��(��[�xK�9�D!E�tt������3��;��q�8�O�4=7�v�,�wɭ=]I�e���J`��$�(�l�b�Ss���};��q�-������G�)����]AQF�nw��9�Շ��G�����ii�e���P_y�ʅ��+������������j��-�酗���#x��F8�Rd���^l*�s8���e�23�����AR_�1!�_�o`��n�7�s��i`�I}��]��g_P��ʍ4c��ر���vO�	=T�'v�(���N���lh�A�[4�[�����|k�9�	e;S�7܃�+~'������i/��'<�b�'�hWQw�C;d���� SW���[ds��G�bPB�!O�hw��O.�񫌟g2
�!~'$��@A�i���@� g���Ԝ9b���R#�����k)�/=u���4��?�0��?������(�/��篭�mI�<:����\+e�D�Fka_*���o@�zD$�ք��J�]�Ӿ�����4|��W��H���<:eԵ��)E���P|_/1���rw�I(mp`)��1\	�0	��Ga�����Fz�bIJ����O�5x�^x_ΆF{[Rz7��
��А�
�ϿH�|���hyςT���~<�'aTuP�������=C�É	o L[��G�:w,���~2#?��)���E�:�G���� �C����ތ�� �@�*��:	<���x�j,e�����B��8.���k� �񃐰�8����-�iI��E��bs����8�	ZN�ns͋ݝ��������AZ���㶾y���� )���qڐR��)[����?�d�$�����}k�n��?U|z�Y�#Q�!%K�wYK�6O�Y�n����z��ǋǟ3��X �>�r�v��L�:�=�Y�PJ���PE��3��é����+?�6:ɰ�\�3X���n�O�>fIաJ��<(J��;l;�Pbc�� d,&���:��U��E���z[�����U�7
��3�)�H�F�~���| 7��/���~��f.��R(�dV���I6��s�y�l�<\��S��"><�������up�������cc���
���f�#�M�;��^�]�Ɓ�[�	�P�نp��D�e5��Mj���R�.ަ���tt�6]���j���T��t�ݫ@�+oO;���p�A7+Hl�;�����R�]k{g�������;LS�4�Aox�e��Yn��-��r�a��t�}Л�?�7R�p؂�H���a�Wg�p��LNg����N]W�E{托`�@�n�ph���6�dAl� P|ck�q��; EX�-�Rx�����o�R�e��2��]��|��@ES�5�G�)���*0tpۂ�[&�x��rb2v�eGܒF�@1%\���X��mec�Pdl���Q�;/2��\��?L�!.��+@$��2�r��ۜ_d�J�wLe� -%_������[���6��F#�7B����1�D��j4,��ӄ�J�tksGJ�a:R�>Q�;c_��IM\�T}[�&ův��)�0���Z|�I.B�2��t�4fL��O�p&��4*�H������n��])�?=�S�����j:���2_N[[�%��K�iE~[
�'��Pt�ȓ;��U�]�]�I��>E�0UB�v���Шt�B#�]�bY�Y][I��k�[�q�`㈫\���첄��6���W5�i(ML���)_��>Qx�Ka?�%�K�V�[��
��0ا�)�[���\ݷ�A+��=`7�������3��E�D@�w��A��� @����_~M���ّ���ҿ�V��E�/q[����­C�T>�sY_ߖ�h���gT��A{}��{&!�":��N#invڟ�<Q'������5���=�ݽݩ���b�� �B�}b%s�z�I�D��9?�S����o���V�U1�R�w��{�q�?<qt��m+ �e������6�s)�G���H㓓�P�=K�Ȩ�S�0��6��=C��,�ܙ��/�5�� ㋗�^"����m��ʧ��0��UW��=�x8+'Q����ҋ�t�����̰1k�]�
��M{v��<d�J+���2/f�3�e?J�����!�p
G��_N�J��gք��\�:}h#�rY��밪)_��AUzw�R|�M�2,�a匙G�mVl��{N��CFx8�wL��aJx������'۹|E��@��&��;��7(C����<���$��ထMx����|�8|	Z ����[�E�u��y\:Wד�Pp�l{[�?�0;7���G��ؠ���S�ϟ?W_v�766�f�'��"x�����/E��b_5�v�Q��JJ�e�V��cΚ���Ff[�1��K6q�բ��3)��ds�ÊYs��qCQ>V�*l���)۪�GF����:(���K�l-8=;5nl���	�ԏ���Һ��M��m���?c���O���>h044$�g�3��f��![j�����KSS�irrJ�O�)<2���b��JOp�o��I! �j�*��xg��3U��O9E׿��3�c�0՟��Q��}�^}(+i�AT>Vb�j�B�z� ��F�U�N���*r~
f��J��&e�5hOS�cުwgq!����)}��l�����I:��-}Gsww�N@�%>���7�a�<���3��$��=���������c.���v<�U�	�RvLc������ ��841I��nP�cŀ����!�O�e�H���{�L�ЛItKJ'Sl�\�@���h`%��q��ľ�ᆱ+��H���ەΙ�u�d���9@Ƭ&���w�Y)1>�Y��� (kz�=�@��ˊn0L�Y:/��$k�O���n�`8�,����z����u'��S�>�4��lA������^"�s��pP�a:��{&Y6��O�I��?刃����@_=C�p�X]�s	?*��[�X�(#_ 䇁Y⡀��M�}�N�wZ����S˵�[����kis���_�������/�ӓ���7�>�Ӧ�?I���)��s>��4}������믞�o�y��>y�6ֶӱ�J�����CgI�3=c��ga'�h<t0'g(�̦{�����̆�c������gk�%�_-3�0����=u(�HI��?�����qZ��^�Y��u�6䶵�l��/�ͣ��)e]J=�f���Q�������8�av�M�Ό}x|����@�\�0��8�r�_���?�T,bP�9�F��� ���6�؝���'^�nn��6x;��W/:�*��l���i �Ǭi ��h���^]����&�QF��	��&�W�!�PѥТز��X�'�e��=Ҹ��'��� ��ޔG����y��Vm˳{��/�'=��.n0d���j�*��?ۑ��$��ݶ�@��r�_ l(����B#:jH��Ôμ�F�����r�٧�O����*��;̷v��������Jz��fY�$��,Y����V6vӪ�+���,��e�K��`|[�C���k�r�M�V�ҋ��B�x�>wU�a_J5�Z;��R��H�N¥��C4V%��::5�g�/+��U�W�)���<��U�ߡp�;?22�f�&������YA��~lL�Y�y�3 q��g,�/,̧���׫����m��~-�"s����G3I�?n�u ��g��.�Z�8��9QF5U�ؕ�^������0�#�@�o3X/)����[�SL��QV>��SL<��~Tx�&�o��=��Wp?��c�',2��{R"����L"9Nn7%u�V=��gH�@�it�
x�rdp�(K�놙�M��(�J"f�I�J������&B��ӏ���}��2��
&*�X�R�.H��'f�#&O�k�́�r��=5<#t��8W#y�����8ߏ�;����pX�f֎��(<h�}��Rx;�T�Pb��ٌ�{zR�4�U�z&��g�׊�L�Sh�ɘ�]0@z��� !�5g=ʣ_80�P^}���j�~�؀�:V�Gp����477�Y۩�q�	�P�V�5�^��m�%AV��<`��Sd��if�w�L �w�<��W����q�w �<F���ؚ�ݷOғ��W/V�YݵU���횄8���B`S��v2{n��B1!P����mix�O4M��|M��w�N���"e��4� ���ig��˷�W�U�ޚ��<k+`F�D<�:V踸�����Xn<�,-�4� G������4i�t-�+%�@�J���m�Q��[�z�����&�]Kܝ���Rz�j��o�:���I��)��ᐗ�פ4���#���S͜Jn�5���$��2�&���ʿ�4������:`� $��Gߐ'��p�t���v�W�8j��r���te�T���pß�s8���w#�?�
�"I�NCæ���ɭġ���r�.����m�ɬ-8��H�=Ԁ���e{+��)e��17�ro|`ލPqn86��_xP��D�β��LƳ�*���Uʭ�a�H&��uj���E� ��-�2�R����ʔ�Vل�ܪ�"�&�(Zo�TWo��zzT��p��hM�����NϞ?K��!��G����t�7~\ȗ�↕cϢ��#Nj�'j�G��j��WV�����L�+�d���j'�UOɆ�K��_z���^|H`s�A�~�;8��/LF?2<:�[e��9��Joe�0�E궧G�G$o:�ڜ�����ff�ٶ��ݑF����T�M&ǆҰ��>��]�ݢ���2 ?�g*+�GG���?I+�{U�����a�&�;������h���yB�`7�����1f@�<c���'����[���$�����8���c47�'������QhoB��Ʋ]"��,Ѐ��T��499�>^��;��
�3�|e����,�f���}��ģ�p�%���� ��a�<��P�+²���&��l�e6�KX�m��e<��'��+��)q��B����[L��s���Ʃ>s�*��D��\��G�m�m��3�ɡr�z�_�U��ff�<�7��y�r��I�a4�YT��fN�zJ�w���؊��Bʝ�! c	������@a0����d�vL��cdxHn,�Hɸ�.|R�SJ�p���L�R9����''����5U��idl�q���r2��S�"i���'�<��&��K��u���:,G|��x����r��2"A4�|�'&�� {l|�8L���ٙY+���qdtȟm�z��Ħ��U)�KK�^6G�Eh?���M�1�1j���b��y��LI�*u�
��w�Q���ā�D{{�<��3�[�{i_��ѡ:���|�����N 8���Um,���s[(Bc�`SӵZ(�CC=��g(�-xkɋ�/�lK������kff_�Hy\J�R�پ���!)�j0 Wu�� �3̬�W$Ne�����T������JC�ph����j�I�S'��I�Vޡ�X��ώT��T_��b��MYXN4�N���w�,oӮڗ�8��A ʵ9�Rn=H���mJ���R+�JTϸ�q�*�#:*U��vm�iTl1E� |��"ܰt�+/����E��ӟ�(v���Pn�V@-8-�1 ��c��3X�M��ܥ�в�xt�.���e�?�y&Wi�(���O1�"�󌭔�\󯰈2�WL�Q��>�~ǽ�l�oB�������v۪N3�[(P�}�������))���	�S��Ȉ�~�>&o�Z��������_r��D(I�L;�W#_c[��`��V���)�^���[Rnz����}�+=R�FG�|uߩY��c���v�t�2�ܨ���
(��ȋ�kɝ����H��M=�q(�ɛ���-	�m=hf2��lC�f��ꃼ�e�~��n)�L(@f��v�V:+��_>5<0@�:���q/,�ץ�r@�S}V(��R��ҘV�Qf�wlmh�n�������2���5�?��O)�A5�6�Skk[޺�܃��L����0恢���l�;?V��0!�Q"`%��n'��m�v��T��Pn��DD,�"��{x�23C��r�?�)1�M�KEi�#o�5��5$Z=!�-A�wՇI�Eΐ��r�Tڴ;�W�[��+U����ԇr���Y�8���4�d��WʭRS�$�gx������;�C.䆞qq)k	��1�w�4���8��ԆPn�9��g�����ƙh��d�LP_���-2�b�~�V�c-�R%7*$3?l�� �z&hn�-��+ ��w�B��4F��p K�лbBD�}KF%��V���=�oߠܾ�HslL���G��ԃ�ݩo��f�������c��Ǐ҃Gӝ{w}��������N���y�[���,3v��!$.���^�Q._4����m|W|`������������tOy-..��1;7��$�~�n�;b�y�0?�p�|��K�f ��ĵ�c	�	�U+d̔R��+3/���]�j�9��������rT��zn2`����=߳keUJ w67KX�sRX��(J�xH#<xJ���^��a��[+'0��x�E���  9C�roV����<y�����Ξ@uR�sf����O�ӧ����/���r�(�gF��%!�Ĕ+�_g-�D..���A�"�U��T&��R��s ��{�}~�u1����NfMؾ½�����wMف��Ԕg��'ؗ�rK�Ԩ�2b�+���"DC(��/��FE��U��W���qǣ�y&ͨo���)|����ޠ㠽ȻRl�Kuo�S�H/�u�x�Op֍m���R��#~+��d����d��fŕw��6+���
7 ��J���~�Ԫ�ݙ@j�+�7eox\�ؒޅ�^F:�
�*O����e��� ���P)��_oۍ�?�*ً����\(G�7�Q��A�x˳�N��+��ɖ�B��a\A?�%���X�� x��8ڵ�u�_���s��w�%�ą�48�gb�~���Iˏ)���!����t�d��~����m�:+N;<k���6+=\)yz�-ۍ�θC����y�1+B�}N�K�ؚ'KT�Oi�!M
w!�T�2���"�|�l=`�z�>�]���(���C�0����d�[V�65�f�-{hG��r�w�H�G�@\�#�}R>���/n��b���j��,��O���AѫI���Օʹ�%�/��	��N)-R�����JuS�"W
�So�p�Ҁ��V�oCo>�wx�}���	�]��H��Y �㤔�ʉ\��/��<��R��?A�a�C�:��y+�]m��Rng��]�rˊ@�����=K)�:܏�b�:��f_�?������+��Xdm�b�ڐn�f�_�K[!�2��8^
);ڪ���vܬXWi�z���L��L��1�E8�K(�����6�܊�[�L��_�[&��������,i�AC��9J(��"E�P.*'���]7z��@8�ˎ�ψS���+�/��8�GԌJ��
�f���H�������-#�7*��w��#M������h��f�v�3�czg6uD�O��_އ��!��h��CP \�^��l���u�AHLx?�0P)l}�@����7���ƥl�� ����ӕ<�_x��߇�ҰFq���j����`�����AZ^e)���
�:�\��2���1?�]�3��{������B��"��u����?
�/���S:%��	O��Ag��gۚP:.%0[��`O�P�� �-q5�}��:m�r�ۑ:�����p]�:$)�����s�u�����QV��e{�Ƕ��~O�����l�6����P��@݈C��L_�+(/t�Q,�=0���M\QwrRS>,���w����?C�K���Pn_�zK�At��R|�[��F�ѠPMK�
flzQ�Fށ�@����uS��P@�7���y;��
j�Q�v��c�Q�;/���͊�l\,&��3��:��
f@����Gbb ��z��28�Tg���)o�5xd��0��"�;��g����A���sr��3���loc�bs�/��&��D���{�F����]�K{�3��+��W�����/5(¡Ēq�bm�0*�'r��"��Ba9&^���"y���|�J��"E���ǔ�v�~�)�R�	[��-���9�DS�<�C�|#�����P7Ж�r�r�/�Qj�:����ٙqH�s���+)��R\���9`vuA�������U)����GVn��\nBQӗ� �Eʣ���E�0�}Gm��S�a���[�\ⳂE�},���~�OHE���42@&�=�9[��A�e۹d�*���>f���\{��{��?��M���XV�L�so��m�@��֬A6򫐏�k��~:������N�[X\��5 y'�V2�m��6Ζ*Q�$��FT���D������`����O�\����7��^�)d	̬�%D�2s�>6f:Ʉ0����3�����8ے2�ecq���Q�n�j��������4)�c���e��B�a\V�T��@ROlS�02���i�cVn5�V�Q�D߉)ۄ�)m�~���D�h �e��5��?� 3�b�0�m���s�Ac�O&�����D��ak(3���{�[�M���.�П0s�������͝��z�3�����묔�fω@������i�
S�2��%4��2sԟ��:�% *C��0�Yy�Σru�~�xzz:����u��tv3k�6��[�]=�rh�t<� Й�ذ; 1[� 7�B2C��`�q�w$���h����B	���Q�k� 7[!Ea����Nj�6�����O�:B�C�P�	^��q��6p��O��@�"ҭ��K��?I����ێ뾿l�-	b��f��Nul����w}qǔ %p��W�b�G7�\��O�c敻,��Y��Z�@�����#7�J!r&��;|� Jmz��ؙhڬ�@�;'f�ٻLC8��ZчCz����������>gG,����g���r%�^\Pn�<[�~c���Т��Ŝ�f�+���G�#�L��o:|�o��OA_����5
�T��n�Y��Oك�@Ly���ؠ��N��r����:ߝt�·����B�B���,]y�O��VJ
�����$6�_�V�t{v}F��#\	]7>V`"��S�JQ� fBF�9���]?"�x����;��֠0jX�-r�d�	̈R�( I�S8)�oߞ)iVy����͍�?(6(3�C�@���QT�:�+���N����n*��3�©4������U_o�Vݪ׸�Y�,�C�H����qE�eV�� ��P�%�JY�����\���|V�+��,y� ��0)�פ��=rg"Y�r[Vݪ����h���6���� ���&�]���������YP��|f�����Wp]��GrNR?�e>68q��������nĵk t��)cd�T8��G�4~�m	?��SZYZO;[�/`�Y���i�����8�v�Pn9#�ml[�Ro�v�%>A}�QМ���WVI�e@�U��n���e�)��i:g��:u�L
4
-�ƛ[[iie�۰�ޒ��(BgRn�	����9p�:Fi�<Wq���+��f�g���\y�x�~p��m8�^�������'��/:>1�ffg�F�ʌ|:LϞ-Iy��l3-�Yǐr�PP]Z��g�J���L`^���P�<#�r]�9���o�sʛiRf6[�JL%��x������"Ōg�	��٦�`�w+�WE�N�ӓ>+24Ч(Ƚ7��++����(F��Y���~��5+������� �x�(q�2#;cR���d���l���G����6�i��?���ʠ(�~&CA(���1���BO~L��r�0fo߯�ҷ5{�M�Q���?������U1ک���@��QH4Lf�@>�a�X�U-�4A� ���\+�Dd�t�A��
4���g�"�p�2`��	yhhXJb�*%>��ud��Y�eK�4>$M��ʾ(N�{	�#�s�^ن�Mikk_��55|��OD��4�T�kFT�"8��Ҿ�HL@%2���>ũ�[�N�2Hc�<�~哼��k^`��@�QMv�2mJ�p��Ʈ�`1����/�cB����. �����s�p��hn��*g��`j:���������"Q(l*<����f_������@��x�ƒ/�684�FGQ9D2*�1���e�	���y\�u����YVa`�.�T���J!����KcApm��O���qV��ǰg:�������=T��gF��L�����LW�oN3����H�}����K�l�`ٯ:]��
 �����b�]ڨ)\�_l׏TC��@UG21��Q �m~��Fl��[^%M�1X.�!�]�+S�f�C	��S�.�K]KM����$:����H�:�NѢ5�����^&''|�c\u1�AL����S�c�vdx���8pD]2K����z}u�8M
C[vZ(�������噷&�轻<�4��^�aWa�gaz�P�˖�� ޳>
�,,M�A2v�c��J�i��(����P�]��[V)Wlc�D����et�G�c����꼲�I�9�x�wD![�U��;�S�t����#-��(�N�8~�sFT��G��d�y�Yyv4����"�m��ۋ�k/�?}�̷���OᓪM�jRpY-���(١/a����{����r�3���1>��ڭu���Q`���T��.=�O�4���<��L3�qu�U*�p�`�`_8q�T��)��+(C�EFI_��>���43���R�|�iT��n�!3��t�׼裸�[8�;��l��\I�̬��"<_��T?��O���1��p�Z~?T���ecK!�3C~���~���]�9��ǎV�X&��9);�J�E[��/�)�45��l��|WM��g���F�u��ۖ&�x���8PF<����e[u|�ʣ�(0Kά<�X%�r{!>U:�.2(�F�mQ��L&�.~�[ӗ?�L@j� �m����r��nצ5���2m3}ES� {�{�I��fo�¿O�E� .���m-�����-�����P8b����\�@/�g���E���b�0?V&ܪT)���V�*@�ϸ�cTLaz�U"@�7���O`DL����O�kۂ�j����y�[iE#UfdYV⓼kb\�����܍��;X�|���+�g,��Cb����Nbu+z|)��L1[#::����5	��:H��8�@��-6���lvX:��{,�c��e���&9��IT6�sh�y�<�Ni�>�&�E����#���h�㡘�l6Q��Bqw�����9C��)m
�0��ƵJ(��iP�����_�b��ٙ�̎OLzo���ҽ{�ӝ�;iaaAB|������� /HI�S�7��m�0�F)<�ǖ�<뤲��C�ol��Rx��DPDX9`y�O��O�wg�Ϭg��V���������NZ��k�އ='�7#�vF�pqH#[�:ʬ�>{�j�f��T^�d\<��!q�hhA�v�8(=m��<"�Den�^� ���p��*E��;AIyX~T��Rw:�I��} �4�V�#3�("��N�0K>2*��O:K��"3�(6$ݩ�Y�xZa������cPʠ�჻��+�lc��Pv��g�[l
Yd�т��+���%̹��Q2Q F��=x�V�e�O�3s8:��֣���<���/�l3ۋ������2�����������r�

7�&{�Ynǘt����PE\�.۝�l��D7PG���EA�y�wl�s]�ϩ�M��D|�#f�겉�
�W�B�^$/ww��g�/)��Ϩ�-�� �7� 엾�����)�Q�ۑ!fn[�O���_�o�J��j_�_���ʸ���#�ֲ��Bْ��]cFV�l���,y\QFѠ7ebՇ�7�\�!��g�'{�Aݧ��}�6�)�ŞuhB2�ظ��,��g5�̊��2`�r�w�^�^�����,�?p(mT����4�f?���>j��p��j�	f��m��}Mh���=����`���N�_�zfE9Ĭ-��AnU� ה�)������M�E�5�;�!GLϰ�x�c5C�l��mCh3��i��Ȏ� �J���N���{%�su��{w4@>%������-��Du�oܬܪ��4��1�נ܂����6��k��Ѯ���"lՒ�E;����6�B-�~�ܶ�G:�u��Wγ�s�[`���A�m�V�s�6B:��ٖ.喋�C�e�6+��L�`�q��C0|(@����0�Ӽ��a2���8P˅��A��ݸq��4��9�R��=��RZW�}��
�zQreKaE�]]�JR7����z���|<`mWn�>�szr�Q��γs▇a���� �����7����ز��6��T�ݧ�Qe\��Y�M	W��u ?p)�qG�����U�P�	HP	%A�	݄���:ƥ"�����IB;��߻��.��߻~�FG��G]F���`����{��R�i,l5�L(�T��e�[(l����C�c����]�s;UƞF��V݊��@�[QQB��O��F��C��D��cJiV'�6��>�ct�c�#=�1�*�����P��1�ߍTm^<p���X�3�\"��WµŁ2����\| T�9e��gn3?�3�)n�/�LQ�9�Tvq�{�s�k[�_��tYq�9D	iP={Y�����Pn���,>3�����D�U�ˌ���D;�\�I��vth��RH�����RIeewgK��S�:on+y��N����҈һ������=�Af���̞���>����e�)J'l�2���'=+���%2H�UY�+>H��lI9e�|��8m~i�iou���aS�`ʏM�Y��xpFYF�n��d���������b��ꕠ�;}�L� �$�ۘ�
qr����d�0����2T�}m�>���A�����_N[����Oi�@�ʭg�}އ���2��A(���ـ��\��F� �A}�%�o��|I}�����;�گ۟�t?!���b^��@Qf���`KӐx�mS��a���/�V^ś@�g�z�$c�K2e��!)DE�e[�+_���f�+�(�C�369)y��z�姟^KY�ʰ��
(~�pPgW�g�x�o<>�TZT۪Ҧ����� \ɥ�x�zj�+S���զҠ0���n�����Ƽ�eb��%��2��*��ß�@~QOU�802���x�@�Y��Jr��8���6�����?"YN�-!���c(�=�Un�ES�t[�|P#L<P�ncѾ�L�Pڍc���/�!o���1���%��󮰄�Qn��?�ܶ�[�� �V��ʭ����J��Q�-$]���d@����JTADk��B���L��8VyJ��6$*�|<����=�^���J��u)�)��W�ymE��X��J��Rʥ�G)�{�tZc��A��J|O�G����. ���=���U����Ѿ[彲�����]=��W�V�Ҳ n+˲��1s��ì�21�˵R��ȕ4�����̭��)$�Nv�Q�4����u�c����x�?�ؿ��Yv%��/7���������<����<���+XҦ���2����˵-��3�my��9�{���W��5):���}(�"�A�j7�@0�d�w��m����s�{M�o�P;����{�O���^��-w,3�ғ�\F馳����-�%fH�$;�;	W�鴵}�^�������Dʭ:O���9���`��DlI w;��q5V�+�a
���@:Y��_�5�r6�S� �DSV|� J,�mR*�W��,�{{��x���{T5�a)�Aw����9)�cа5���sw��B0??�%��~)0�^�e���ʒa����+�\��ܑ�˵;�zA���ͤ��I���O�"u4Jgsk�a�'�->�l1�ԫ?�r��� ��g��B� 33?]\�EG:5�j����ue��-���[~���*�E)��ޢCw�3ɍs5J��v���(����7x:�E�v��c+�����O~�s�?�	���Ga�g�}�2�gp!��DXȊ 󢜑,(샆����r˗�F�����@�:a���w�.�>z�~��G^�������Gw}·><��<=T��SO�{��[NO�}��E�i��3�Uh@�.U�X����{w�ˬ�,�#V�q� �9߰�pG��Aۢ����Ϥ���!)��=����#�������>�Yjnn��/�}pX2�S2�9mm�����%�%�$��$�J����v�(W,^�_�W�.e�;�W��ƖR�"~�n�O��"��5�u�r֐߉���W��BX/����N;2hE���7��)��<��wM�V&�c� Tm�vʪ��[�,ߖ�2:�!�����oG��T���r�O����&ܮdr��g'��,�c��r�Y��;�9��_D~�D�Θ;M���"�8޼Nb�E��(����O���:�:aB�r������
��[�%��?+�'(��w!cX�V��s�����a0zu��ѲP)�\���:���xd�����{@�ƬmT<�B�oht̐r�������W�؇p}w���i~��6~'��w�x�RL���{*Q�-�����4��(p'L,;�Z�D���S�uȅ�܉�˧}�J��Z)�=���_ >�r�K��W����pz�2�Ҟ2A��-ƴ��4�Jʤ���cLU�"D�(��u�_�p"�ȑgse�M6�*\���,�����<�g9�S�zC�cv�C�q�#u	�4Mi0�P���h0��gϳ�|M�����詊.-"�P�Pp��C�b�g~a��J��b��@DB)�+��b3x?n2�Ua��}�\trz-^�Lk���.j_|�!��}�/:'�#�x���r)SQ�a�%�C�A(S���Xb� ��F��Rܜ�����[�G�B�ç(T(��`!piT�زP��;
K�����Ã���Ŗ��K͡�rM_Y���:8�A�$?VX�����^jFI�F�E�=�g�e]ͮ�ű ���Idw;���ꪕa�o'�����E+�SF��OK_&��?.\�\x�+܇|x�ge��	\1�!
x�������X�:�������T����s�:
q7����dkJ�uڠ܊��e�C�A톊�z��?�DDYюX]%��O"��22�*<8�6�)m�}�H�	D~�b@�`�,���r���!�Ŗ�M���-��ϩ3sS�:��K��L<�f0ŁVn�a[	�R�%ǸǛ�g|��Q��2e����
?oCр���k�{<=zt�+?3�ʋ|���Q�9��L>�'�]�܋���<K��N�#Ck�Sge���Ս�`�y�kx�%m�mK�/����|꿅K���fK#h\r�3`0�=�JW���Zk���{���FddUu��_��{��8~����z�V�i�|�&Z��.�Y����r����ƍk���l���V��]�b�pj�T�R�#����>H��̒�c�

3��2ˤ�l�4E�i����VLy���'��ۇ�s6��'��;�'�cE�mm��T�+|I���#Q�/#�(�bA���%��f���ůN�)�8�3M��x�k�YFdWA��X�p�e	ߥܾi�6�>~r�7d�3U�^7Q�"��M��W�)P�g�CC��H�rۣ|qbB�E�=�$�����rK��%�%[$F��ǳ+}a Ъ�U��V�K�&��/g*� ���n. 2-4=�ψ(���@6��c�(Ћ���B1mܡ
ʵ� g��
��8 �jH8RiPσr�`kC�3t�V��2A��4�v1��|�=pR��'A�1+�l�-#�g'RHT��ِtDϐQ]
���
<�[�S��Mp~^h�&�P�H�eόbhT��f��.$�W�����A��z���q��w{	�ЛN���{���{���l\����rz�l%=~��?_IO_��g/7ғ�k�ɋ��bf+���6��I(g�����ߙW,a�[
��w$��f�#YΚ�	�%^��J�:;vH�\��'\��ս���Xv�ю�����y�V7�G�O�v�6���֎���s��徼����Ӣ��Lx�X�z6F4*�� �%�tQ���68�W�h��Q~};�� �X�������8����Y�!�T� �
�1����pq��Rhyofč)eFjc�T@��"
1|�$]7�cB;n
c$ N�ؓr�Y��-�����S��������K��V���C�e��򺻫�P�Q�T��C)����pF��h y>p�ʇ���=>ܓ�+����pR�&�e!�A�,Q a/��c�=L���p?�ß
�]�6��k��[��ܚP�@����B~}�̄�����TӲ �C����E��<���h�çw6��H�/:�ς��D�0e\߾Ø�(s�����ԓ�K�h3�ݺ@'�����By�.��Ju`�&�ӄ��i)��q��O�K��B<�Z�A)�=N36�Q�H'���5,�-d7W�s�5����4���w���:m�;z�w*=xp+=zx'����������0����p��3��e�S�*Y���Q�99I�e�Fa�������={��<y鵶���3���ҥ�i�Y�g���Ϟ���������$���?���r�Q}Q������V��<S�*S��K�CCSʒ���6��ϛ|���]�+��mld�Qy#��1u��ϳ��r\�b�-?b�%�3�n|i��k=�?Θ�J��W��b��2?������i�J=u�3}�q�ǛL�~#�����������K�0ᖨ=� 8�9z-�@��09����+n��b.~�I
�@�.gR&P�AXe��Ư��C�#l8رfh�bC�bD!�/���F4�z�e$L-"X��=h�N9M�G4�m|������g�WB���13�d� _�븃�LvE��Q���nr��H��^���#}�&}�7�P��=�8�k��x�=�
�*@p����W��U1!����g��=�����2�]��<��=�޵*�r�W]nKaܳ�M�+[iuu'-��y)/M��Y�����/a�w�P"�"[h+�˝H[�Cit�0�?�?k��t*%J��-v�r��pN�C�y��lލ�pd�7	qC~�~a#�ί��9�+fw�")���|oe@���XQ<�S�駺��XL�@]Ԏ����Ř �zD�x� +߅&����Vz�r��Q���8������B�W4-�����
P�,���)Ť��3q��b����:,3VNY*@�b�ld�vy�M�� ��H'�6����FZ[Y����ںG^��K8!����i޷�1z�,�X�����%|zLs�f���l0,E������1"]6+���
o��W<�I�r	�RK<K��&�z�4���sz���<;.�ì��IlR°� ��^����r�F[o�arYf뻌����y\ �\�]���u�EF˶�l��m�%\.�r�2Q��9�Wӓ2�T6�ť�kq�����t�?��'�3pV7K����D�s�e3ò���=��`9 ���DT�S�+!t���Vn�i�H�вG����^g�����/J#8qz8�ٙ5�m��$`��F�x�w�*^Jppp.y�VVԱ�YomH���;u�[u�eg��{�G�2�ȆU� ���p�3a̒�i����뒕��/#>$���= t\(�(�(�C�l�)��a�9>�����e�d�7���P�ȧ�U� dn��?�ǝ�p�����L�(��e	,+b��[�^��,�3���eC�G���dI#���Ȝ�&��ȭ @�:�

��?�ǺD��_6��ס�S�o����lA��A�ߠ��!�\B�7�U�Ie)]��ƚ[fOXsk�_�8��Vu>d���S8���//���Y�կ~�|5����0*��
���%�����������IlW.�/ְD@���Ƹ��׈�_NC�l�[��L6�qF�܀����x�o%�Q�F0���n��SN4
W�.#�U�����n��4ɇR��S8�8ȍ`�� %��Fcc����$�lH��0��n���C�x���jT��~��_3
t]`Lc���u&�	�云X���8���H9�ܰ�B�@Lkf�԰a� �Q�4<�2�b�r�&�GN)�̋���əG��J)E�3A%s'A�!�ChgzX`%�>R��Pl�Ti;=�i%|䍆����Q|��4��ӪrDY�.~��0��������#���:��2����a.��qn慯qds�e�!�E������n�ʔ
���|����;�Y�����4���a���(�h�@y7�.��1r���z���輳��v���8��<��uʖ�;�g6��9���(/(��k���iU�顔[��p�����Lw��e)��j�zv�30�ˆ?6.B���%)��q�aŕ��#�'�Zq\Ԛ�S������k��g���B�Q���Y�Y���>�'-��i����K�����ȁr���y�YG�����x𙘘��a�������y�a��͌�ql�TZO�#3}�L;�^]Vr`/�b��߳h��� ���q]��\��VtPȤ���� 2�|A�P�^SOݲ죚�˰�g�[�v��1�)n���9�K4��s�e�#���ݛ���[����4�Y�]Æ<��bYt;:���7P��"��!V�̬��'Og�_=N��ç�����02�t�����$�@d?6*�7�cY���?����+��Ǡi��� ��9p4��G=s�)��#)�ۇinf9}������4;��+�;:�T�܁W}!f0���DP���v���7S�$�{�y��$yTd���K�=���Αۨ�[��̏��ϟ���/�s6�[6�?�;�nD��ʨ�HE~�g=P&(���9��N�Ed�;'
��+,�Lq`F��d{��p+�w���N?��{��ß�;���&�qs�� �M���w����rz���d�a�<�O�7o�v�Ԟ:k+��Oۻ;����xxM����[�Ey�<.�ȁ#�E;�2��G�8,ӡ��"�xd��%����ٝ@�i�������?N��Xj��6eK&���$�b���|�q���y�����Ӧ�����˯����o}�]��.�e #�K�<���GH�䙌�ix���E5�g�9�T<�gn؅(�0ma��|s�c�� q�
� �
��%x�P6� |�x6&.8����>��{*�����I��x(�D|!������u\���WF�Xl�p����+oſ�ɥ�O��8Cs�#\q�q@9"0>�ġ� Q^��*Qؔ4�5�K�F��bE���+�/����w�&��c�'�4eI9
a.�z&���J��*��<U��QQ�ܘJ�;G��
��!�TIU���� ů0�P��-ߩ��d^�7
��L���!�D���S��'����iX¹aS�(�}"��,�s� ��`�%�[�?#Ԭ���RR�𨁈�N����R,!�,!�(��(������O�mA�w��('���'�����<ۼCwd�}��q\i�~x
��rˆ<:�\�@�Ά��u)�+�ien!����&��%"��(���"HC� ���V�]Q|{�9&Iʜh�X������^�͈
��� n��������ϊ%x�D���k�1�1�d��A��j��c�sZ�|��_
02�lLc�.�hT��f6]�*m®o�;_�G��CL�C{�2���ƀ��g���V�W�ضK���R��6o�u�R|X��H	�<j��eS�;�q�[I��Op3�<?ӹ�N��!ߌNBW�`�o4pЌv��x�a�{�{ٯ����s(��������l,�86n��<c��<
��[��h�8 ��ևs��Iw�u���H,���C���󴹽��Ĉ�#O�O�;��m9�����',c�C56:*�N5�R��ׄ]����C�P}0�ȯ���@�<>:M��iuy=;ZHK����I�p�
��8� !(gu���GA�R(d�� l��G>�IB��!qc����>�Z^��a�R(�$��mQ��'S�m�2V4��w��O�x�+��K�ć.[�9}��zv�
E����rG�i:zd���-ʣ�ZVnϏ��`_{z����Ï�I��?���Ng*��\�tGx0�v���3��X���HS(���o�5u��-���6�h<H_+��C�T5�^Y1uG<U����k�K��I�*���[��1�D��u^a�qN){�B�=��	�it�vă'�[������Ԏr�K>�{d������/���Y������zm��TŤ��IO1ʨ�B�,��}b������ f *8g�q�V4:4�ܠE��I��q��D�P�P6#�0$T �Q%�R�ԌQ'�P9l[�Qq����g�d
����sz�V6��b,��vƫ���#�.=y�����KHa;^�PL�@��m�^)�6��=����y�������/�J���4�A�n�9�l���_1_h��q�8e�G܉�竦�T��0�Et����F9d�卲<U�����gQ�=�!A�r����u�A ��^�0�0vfҐD%�OTzlx�x�r+npd��/�S�'�wo�����	�sT܁�6=Z�k�G��=r��>�Ru�BX#	Bh�*k=o�[_ˬ�Vn�A��[�_F��	� �O�w�1z��d��{ x�4�نfVf�v�=	4n���|�:m���΅�)�7��1�:�=���A�v�����'��y=uKaD��*��yHe(���o(F(��I\�(�Lo���ֻ�"%>��V8��6f�By�l�����FF%�G��3-K�D%ꝅ|L�6iq��G�D�;e.��;�ŝM(�� E��n��6��.?l2��H���7�Ti���-F��3�(@*���K�9ۮ��kS�s��������H԰�R.�+J�s}�@h�&�)���&(}3��r�0|�H�|U�u��n&¾l"=x3;\1���5xlW=cC_��
FLU9�2Q����f1���J.J$,�t�����J�T~�pp�d�t�	���K��rˬ$�E�(������H]�t�7D~�A�[ώd �� =�$� 4�r����)�{�M�,k������'�E����+B}����}u�rk��'ɿ��:i䉕[A 8=���N�6��ڧK���g��V���b���t���u��2���������<M}ćoTn��rW|�}�vg/�2r��v�rˉ=l�rۣx.)�O����GQn���[�ݶ�˲��rKH��hA�(�[��q��n�6i"7
���9��u4��{�%��x��������dGgUԴ�m(���Vn���(�mk:�{^Snŏ��n���˿~v���O����_�����^?r�Ϙ����BO��A�ޮXm!�S�1��Lzʘ���R�� E((]�zK�Ő(�C��c�(Vn��p���K�m
8�B���1��!�Wb&~r�)P�Kz�;��V	�-xGC��s��Ŷ\rx��^%�64���ӂ��|��|a
=B�
!nQ6V�f�U��-��H�_2�*�W�Ӻl
�\)&�#]��?��2$����W�!�1��T�Ε/G@�g�F~��T���*=p��Ѐ�.�%#u� �#��*窬d�ʅ�%}E�䄷#�L�#�(�v)c�3t��t��ʦGKYZy�q�"�r��U��CpN)������~͌�G�����`�T�^u}S����-<@L5�x�?�a����@�]�<�m�T�%�LLz��9�>��PV�r+�6�$��Ζ44��c?��]��]_]JO��*��o�]Z]Z򹝌\�z�쉓0�o�pV�dP��dP��Q4���F6��+Ń	!�e�E��	5�G��h�ȗa(����j&ˤ
:��N�e���쪾�7厜��%i��FPfh��p�C=/i򝺏!?�� �S6�'�ɔyG7�L�QP7��r���޾�R���M�3�OA[�l��I^�����gʛ�&ldz�^W�[pogiD��~nձC��oc��ԿdH�!��&\֊�r:9��A�W�|e���X�"�6���-k��x�щa9��5�)Cl�v>g)�Xd�Ax�1�o\�u���/�P����m��������g���z&y#��g��
��
�ʄ tT�?�?��Ztn��*m�V���3�"�A��Ҧ�D��_�9�F�`ӆ��Y�U�iwX)_ �NdF|�r�_Q�]��X�K��3�Ȧ�c�G� 9�ȋ~��RF�O"�I�����E�u}B��ys����w}�@������V�mKLK�}7��/>NwPn�O���j�H�o��@��RVn�r;qI�][^�r���c�<�)(�ȓPnA?����?�����T��M��=��L ��6�9����5���)�k�@��n��Uʭ�%��P|u��-�f$��`�o`cm+5�����/�����^zyJމc�@�M���(@���"9T���*���h�$�"����"SQ`ҧ�. �D.��l����g�S�h��W�HrG	­T"!�Q���[�U�4F�a\9��F�i���+'�o<�R�1r�����.%\��4��p��\��G0vT���U�Ʒ:��i�����S��-?��t-�N���Ttxs y49�w��6���ƺ֮n5Ԃ�._�؎[w���vO�3ǹ������(�����0oW�h����q�w�����`�;r�3G:�N���t:4&n��yz��Ga<��yA�7�pi�lo�4>l�~9���2�?�@��Y1TU4�� ��?4�=�4�,\���/I7�"���F;&� ��<����+r9\�Ν����)�s�W��iow[�-� �����{�g�)��+Ҷ��v4���4�tgD?���1�@F�|yӐ~�qp�md;oȻ�7l2?�L��L�1RKX�X�#;E/�$^X^�u�
ENKvS�P:��ZOC�4D��x���ǻ��/��V842l��;6upt����=NbP#��ʏ2\6�;����TG����:�/q��i��D���_�4�"W5�=?c("��A:��:���T����jlܠZ�7����[��T��,X���-֨
_H+~QeP�zD�W�3!7� �uW�P��Tr�tM5�J�eI����aȈ��=���:�Cu�9ǘ��jw��9���y�q�\��-#��Uy6$��Ȳ��_�Ë�@��WuC����w�4إ�V�p	���AH�6�|��*g?��0<_o�pw��n�q���G�-�r��d:�{�	Dd��`�Љ�ߑ�{s�7gݲ���_��`UK�r�^�tʲ"�A��z������1e�N(K�����BiD^J��J�_�=d$ax/y���!�D��bJ=�v�xh�eC�������jʘqCN��N��#�m��\��y� M��%c���.��a2rU����(@�k0��P��_���y�3�y���:��~�Y�9�.LӵT*<S��Ķ���,�v��ΊӉp@�o�5��((W� �B��U�bj���܀2���gw�#f��[��8���q�d;����*"F�
���hs)X��u�'˳��6W�\y���Exg���8V�Fc��#�ԛ�TYb�� ��nL�RB:�ȢL�%�AoZ�y��`�t����0d�D<���X�>b�uLo�� �~k�o6���m���\U������'�)�
Z�E�̓�;p�}`�/�#p��n�@��o4
//��ӯC��B�<#��;�}�:���LͶzͭD���)�c(rV����ѩ`�AtB����2��.O葕]+�Q�\	��V�S�_�t��3|�٪hNv#����3&��ݞ�,2T���Q�mEN�rͲ2�[i|�,	���Є{4 �e�!��h�ey(���[��ah��{��h��EN��;: �1��"� ��fG�&�ؘ6�]kL�����*��}U��ʅ4��Ȍ�_q�@�� q����<�=n-�D
���ۦvK��F4�!�@�&����K���\�R8ɐ���x,	`���|t�j��鯰�#��Y�$%�;�˗^d8����a|���Oস�u���(� �ijf�����$��25oR�/���r�2��^3�������֟�'p��qڋ�eدs��`��I�dp�7��R]��u���X�T|Rҗ��M��W��¹8W��+��Pfx)�vJ޳U�aj�?�]�1t~
�aLn���v8�Op�� 2�rb��b�u���xɀT WP4�@��ʱ!���>;*��+F���-���Q��j��H"Cz̦"v�����M� �����%��&�FS�q�����;ᔘ3�X��9�.\�?FI#$%a�e� 
1��u`����:�<`g�`�"2r�D/}�`�2)��7fȟ+��&" 3���rS|/��Q��60~����+�K|Y����]��S�1:��SFwX����/�]z ��A� g�r��G�����E+=3��;�Y�"ʞA�s��X��G�1��iT��6��rW8�w�A�&����T�2_��� �xq<$�ʭ�G�O9s�l{�r��/u��3�I���e����8��\��H<LW��Y|���7�=��u�QJR�%RT���Ъ��ct��^��D�П�	 -���[�]���n��ad>v�ӑ.yFd6�k���O1���76���U:%�VFF�x.<˻G<##����G�o,7�x1�J��#��!��Rڬ��	p �(��A^�y��Q�{y�_��K�'w��<�!�1��e�����]���n$nk�����a�OF�b�����5��4�Onq��h�|��\�r�7�Ř#M� \���E�_�7�GL���=�[��)�d��;�l�c=r�{�̚tvs�A��Yf�
�՞:Y�,������٢n�;�I��	�DQ^Ś�Ɏ:�=�V���,36t|�|����3����2�̆1�wv�
���t��}Ї:jd@G��(�����Z���Qvc`*�o���y�/�<cr��}���)S�+�������m���o0��w�)&� o��+n%J�Y޻�π &�z4�\����f�T�Q�ldyQx���5�C�s������Q�0��5��F���X�d��{�aD3�N��!���*��������f�7����,\�C���V�X9��&	�!fþ�����c�S1�A!1�K���S�NлEi��8��˿`������#'d
��@<��Ts��,M3�P^N9NB ��D�U�(�� 7H=3�z2�Jk�p"�l�� gD�
d��pRe�P\^W��ש�5�pȺ�f(�x�ل��"=�
#)m+��4s�$���X�f��DW��Вt�Ҍm#]�����G�Jd��|p4���(�*�L��0縌�h�H��F'��Cݠ},�Wc-�����Qg�0���n��e����ٱ;���	�QfQp]$����[�{,w���������z��i)¡[	�߽<C���2 �i��I=�<��(�LJ��P5$���妸�}�l<�p��i�n�]O+���d��|�d�t6�P�.���_����:l�kQ���.`� z���X'�0�f)���a.t�3�)�,� a��x�^�'P���n��&dF-�
��8���q�������v]�/�G~qsx�)���݃�9�ղ�Z���W<6�X����)t�CބL��d�x+x�*k�yȯ5��G�cJYF:$m�;nQ�A�ƈ��Z�O�ھb�~��
� 9��҆.�L� ���/�o���8P\��Bwʊ�Q����Ph	�� _P�d>L�K�X����-� m��D�<�����9:>a�J7��K���)�M0�>���k���m��$�?���`�(�y�r�f"�2�[����_���&7�}�=_j2����:Xg@&G���-Q~�,�!�Z|Pxʵ�㋺����BY>���p���g�D#�a��0�Sxǐ�n�d�D�m�҃�[�mS/��+��$�h�����h�n�ثL�K�+C<�F����(�-K��������Vz���f�*���(@�&����P�E���%L�����T�vU6���D��;�	 ŀ�+#.�@����VZ@�|Tr�


�B+�5�RT#�j�7����M7< ���P#��2�e\�S�P�۠�>
Gy��3?{��eÒ�)�J�p�h��<K  q,�r/L�?�H� E+���-�����E����΋�s�A�~�t�7�(wRb���>G���VhE��ظE<x��FV���2^||��ﲲ��	����K�ʙ�b�w�P���<j�GI�W��/�H��S��5�\���	�1���	��E�/����vO^��B���rw��4�<��u��g �<�7�w�W<����f���p*�(R���h ]�2(v��n!hOV��| yu*J��@�s��+%U�5�.�M�D�KG�;��4�v��~����R�'ٵ���;������/zz*�0���_�~���Y�zt��ëzB�E����R�7ӏ<��y�|b��P��1Ʈ��O^ʖ8p�[��_�I�vX�/ܲ���Eߪ�"r��V�7�Z҈�%bV��v�nt���
���h�c``DS2G��HZ���]#?�I�EW�ڹ��P>(����hŝz�g�Ǐd�;	��e�` ���%(�� �c�*��Ӡ�K�.?Vڐ��d	G���͝"!�`�ȿ�M�즮�?�~}%��/&>��x�-M��)�gA�B	Z��Ǵl�� h'Py��Z��;�Y���0 J��z�s|�0�;y�M^�9����\����@\%2?�w,����5l������ҵ������S!�������Y�4���������D�?��?҅��F��~Wx���v�s�~���8vn�c�&FS_wbU���࠲#�p�17%��c Y����%;ā���c���#z�����&�����;�e�y��߱���ȯ��O�Y���K#H�H/�Ǹ~(.�?���G���q�l�<D�g�����^s��(�8ш�S#gFw�F.̀�F�dRP��{�6�i�)|g�x�,�d<�T�T������uPv)0�2�#bU\��(D�� (� ��2�|��J�<C�=R�u�jIv��(&�3cW����шMz���`����!�Q�\Y�vP��T!<�J� 6^��P����۔�Y�Uy��[���c�ۙ����M�Nb`Q@�e���.�L?!�4B�d��7=�rpm��A���&��W�s8>�a���րH�0�Qa�w�����\�   3�D��#F�U�Tϐ�TT7 "h(��@�5]$�?⒛���<������Ql���l��)ad�������B-@XB
��(4>x,��;h���AR��?�3�
�� \������ ��v�2�_���ܴ��g<c��ϥ���lx�|����F�ȶ닄>���6�nn�l�6I��H�B��������i���3�Qv(�P�PT���ˊ-�Q`�t�<���SɄ�3��| �_@Y�VLί��Q�s����w�~��!ԧV�G�'���1�E	���qQ�,�� �C+	+DYF�k_�����nv�������;P����P�J=� Cf�!�Ƨ��{&��Q@F���|��P ��ٿ<��X;_�~\������k�U����8*����+���F�qP�a��5�Ϥq��:�oU{C8<ɋ�˰Q#d��2v�g|�3�`��?�N^KDG�;��rD+�Q��>�����_�{	��&C��h���g���{Ø>�9e�,�ئ9eY�p@���"��p��w���Eٿy�4��,�	���μ���\Jz��2�(�@z*��wq��Qv���0[0\�7��V{��#y���Hqwp/ad��D�En�v��s����Th��bf����3�Q��9i�b�X�.�ȸ@/���h��|����D��Q�zqax�_ͭ��S��^� ٍ���33AA&C�q;�@���+�O
�x����4�Dz��P\�Uɸk^����OV�D�^ح���6o����Z2�i�!�?�o�a���$_���%s�JΣ�J��5��_(��4
�-�ڕng��K8t����������[r��T���lW��ڂ2C�ӓ�H����{L��R"+^�%�\+��ɠ�Y
��q�b�>�g���O0� A�;��������U��N�E���"�
(P�����}�t�=�I+1�
g��e �5�v8���H�O(�Л�m�E3G��Ѥ��n��TV0W���+#�xu�l%��Y�<4�
/���:�b��­J�or7�e�v��?_1�:���$�у XP�] �"=��c��b���I7oN�[7��`�y�v}u-������u��\6e��x�h�r�	Z=2]���8\��cv���	,��{-�?�H�?�Q�U]���3UKv�evd'������L�;[�#�pS���N�PN��PśԿ�S����(e��_@��c�[%��2"�h�e?���x��X��W^ِ���xnȤ�}���/�k�⠺�_���檁w�����q����IIs+ju�&J��c�~dI��#��p^�7��?�o٫�Ku�v�>V`��lVl+嵄�7*�����	��*l�ϵnQK��IK�r�^�γ2�?�i���ѱ�aec9�����>;9��7�t�2V�,�r
�\�Iyj��hg��#��K�1�|-���+m7�s)�/�i֗�9�R�x%�Ð_��A�0~��e+`W��[���S��2��e���^���*ۡĢ�1���1pZ F�c4<ܲMa)��+C}��m��Ѷ���(8:��� {�[΋ھ���Ͼx��������	� 5�4�VV��B�y�@�pp�EQQy��G���T@H*��a*ܕSN����NsF����h�΄���
e��
����o��KbNA��d�R+e��]B��8�X��h3�`K�@D!w�if�(J��,>f唑�"�>R�C��
Oܡ\EC)�����vG�)@�.C�϶����!�[1
�S�h&�O�Gio�<��X㥸c�A�݂�]7󊾁c.�k���O&��U~ح+���w�+��/�!4�Ti�)�
6�ݛC�S�ο~� !���0ҿ����D�č=,G0�\�#O�Y�r�9��'���
���(n.o*7���-��K �Уm5�^����7���r\����B�S5@�bD(��\�z���a9ȝ�63�%�cYy�4��N��1:F�M��5S�ڎ�2[/O��,��i����`_i+}N>`�$�}	����ۖ����?����V�Me�!y±/+�+iyi)-..������D�^w����������<;.~Е(^�>�����M�p��_7ƌ�+C�+����O9_Ŕ�ט+1���e9A��{�4�5r����G�����>���P����=nh;��!::n��!�)hC-E�
��!�%w��&+�
V�h���V����X�>]˻�����������⍦��ݰ����
��/��m'	(�#y�C�
{�e79�l����w@d%�J���#�E�Qh,A.��qc|%�H�8"R�q�&��IYCC_&s��=�\	����9�!|��x������$�����e������_��k������G�ԋhS%w�IJev|�βd/&xJ4�M�X^��B�$K��m�+���䱗4"7%�ɿ;j��g�Da�U��d�d\�+��]���Hy>�I=]�ijj(���n��O?Lߺ���Ro�c��9��`� -/,�Ǐ����426��}�ô�������V$���C���|�T���T�!_�2�}��d:�'���랟d��w=s|�F�&�z�[��` �d���Q,�]�L#�ilrR�t�������\Pߺ:��!�F[��iJ{���l��󯞥���#����C�Pa���`c��X�z��=m�+�GE��/��\a���H(�(��gݖ�9R!�0D 3�����ꇙb���^�)�穿�#�w���^�Y���L��CƉC��zݜmE%�ނ�ʽ�5���r��=mcc'-�����]5�(�R��]ڌbt)4	DQlOE)۪<:?6:�ˇ��s�39]!�KEb�����0�3+ꙛ��b�=)���iiy7�����<Lփ)^{�"���A�+<C�(���{�9#q�D����Ke+anx+q�}�?��������#����\���p�{�������i�2���|�_[I<\+�JǍ+2J��*�!#��P*Q�Jx���*��тF���xΕr��Gf7#��r"	I�����4d+�ƷJ��7g���J�����c�:U��r��Xz3ۿ�r[�Y���r�����J��H�A(�,ݹ8�"�]Տ�4==�n�O��N�>w����_r����fgg������׀z'�5�m�.��2�5��H���0���q)�|��4��^
����0u>��.�o> J�]���b�d.{���Yy`ʟC�q�Ԁ���4>1�&�����[���1S�[{i~a%��	f�Ո)<'�C�B�R��{�?H�nP��o�x,�c��,� >���c:r�|��K&���.��Tx5�8~��t���A>�O��kɑ5x&l�����Ɵ�#�%M�I�K�W}���+|���� [4�0�V�D¨�����k�[ŧ�&=�Ox�#�Y��W���[v����XdR��r���D���s�wܑYѶ�`��?��	�o�.>�%͚~b���_Un�%p��((b12���a|n����Xd%<Cz֋dL�����r+yw~���;o�	)�o?��>��G�m)�é�'����N�����n({������X�����-)��喣.c0�+_z C(��u������A��n���(@~��Ŷ{�}��(��4��~������oUn'��v��R'�`_�_ʭ�v���&Ŷ��Czd������U_����7��9e�/���m�EcY�0�}؞&���s���'If��FMQRi=u���r˴*���QۼA=M�$��B��K^'7�"��ґ���8���Q�grX�h�us"�I�dJ��
cÄpC��s�`%]�(Hz4Y�:�����aZ[ے_TO�����T���>5�,t�@A��!���hzft�XF02<��ޙVc=�nNO����Ԏ"���g�sI8�(�8�?��(��Rnw�O���nz�tY̺�ܱ�H����͔I�~
%S��C�KP�)1��f�58"��C`D!Xx��K�|�g��T&0�;6�`(}�����G�vYՌ>!����j��-��@�y�rKE���
��)����Ih�W�r��黕X���$h��� ��-���2�!h}�1h���*S��:.+��M�b��'ҰU��m�Tz�i�:%嶥C��S�)��ʭ��OPn�j�[T�P|��+�d@�k9�[(-ʣ�~*>�8!!>=�vU?��[n�G����y�a���������ffӳ�����Bڒ ���[�i���5c'J�7�^\����]i�N�k�k�-��;*s������	�j�^�$;|G#�N�\n�6<:�n߹��ݿ��z�VF��U��o�4|������+�K~l��J.]Q@K�֋y^���7�'<ˣJ%�)y��Ge�p N^������t��U#Z^�,�`�dg>��$����r�1ᔿ�r��U���#.J���N��!�\pD�8n�߃���C$�#��%;ԙ��ptn�q�%��۸�C��T�ǖ!p���p>�n6|P�}��m����k��FnvqF��h[�Gg2��@%ʾ
x2�G&@e:-�g�.�ܒ,��x�qaB(����M���G���=@,B-���" ��Vz���^��[��M��B��0����45=�{}m:r�=L�l���gϞ�r;:$�[��v�	C�2�/3��n��z���7z��+�Y_q~�,϶�����[�5�'N�����\�%N�%�!ev�vlD��q�ܲL�%�{{`������K���aF}ow?5������/�|���z�;��Z�P�f8%+���M���� ތ������ۏc�
kZN��=���2�Rk]8� *x�V8�	����� >gc�`�|.��P�m��{w� �u/ݿw;ݒ95>"�L�C�R0����@eul(��������`��ʹ 
2#o����\�b��=J�z�,��IEvQ��bk�Y��Gz��N�����]�xS�8*�wDx}��dX8�Vc>$���@�Ï�)�idDߕ���A	��s���]�\���~(���63#��d�;`���_�SV��Q9J|��vy.���z:$ #���d��m�Rk ~����-kN��������˅���ύ��Q���#��E���)k�b�ܩf�Jt�K���������s�I�A����M�C�-����.ܽ$I���s� mA. o�%���섷�;=�%��_3Q��k�y��퇿pԣ~JE�B-�9P�PCt*�2�2;�0ku���O�Ug�%����Y퀜��Wwvv�&�ks9�2���ϓ�������]6'Gwn��M��qռ�ƻ [W��M�Q,⯥#V���|.�� e�gd�ºa�M�*�^iԺ�:%����T�u{�rkLr���S��=��.%weu=�3%��Ý9FnQV)k�uDOJ��E%�v�x���xJ�ʭ��Cs�I<�l�ĥ���q9a_��`4�5�-˝l�ғ���,�	�8��C�?�I=������	8�l�#��>.�1���F��5���C(�Qμ�W20����������N��ӂO6�?� �3N��(�o�0<�Ǟ0%/���Q��/oUD�鍀y�;qRF���O6iK�Y�U_�{T�{}my_Ow���J}}]�@�xF�C���M���W�ͬoO�b�Ma}�˝��@gW�ŭG�{{9� ����M�љ�6�v��� :�yjV��.d������q�(}����Њx����-)r��vvw�&/�� exw/mmm�#�k>�]'��W���N(���te"������,J.v���|Q�WƸZU:�Qϐ�>-AJ.4h�<aI_9)����N�8��s�`�4������ť������w�詗�ԩz�6����)!'n,P����A�k5Hy�� �q�g����^1SwOG���4c���]>Ƣ���8a���j&�"灈dB��#%�Fӱ�C��x�sk*ݿ{[�㸔¾ԣ�ocC��CϭU�k:�}�'8��76h�n�\Izla#D�����VZZZNb(���>3P82f	@�P�2��h����LJ�F�F�����:�r�kpn2N�㢊���^�K)tFfON����`?m�o��kY�2����9?�ih6�wp��M)�3*Dĕ���7�5��.� �)kW|�����+�휏l��V����j��w�ƙ:Ky�u;�r�J�z��vܴā�\`0�Y�)�M8�#l�v�70���+]g��/4�����UC���zp6.�w$�I:ldp�Q��ڄGn�jec#6~��A~9T�t0-H4c5*�<��V��/�i/�mY�sń��/6�^�=�Ad� @�!) ��iۏ�AG��ɩ�[)��L���e�r;8أFF2Eu����f�L��,ź����f�� ���m)���>39 �x���,p.�`�^u��F�����x^�rա�������l��4��g�+�WU.�1:��74����)j���ّ\^^�R�����a�U :;%�s�+6����=j(\id��1�
n4ā�����o���C�i����P�ilB���,w�!� �%��k(��k�S�݀L��P>�y	�÷����'��&Г�td��2����q�Y`7�G:��F+����*��FTw��Yq��PO�O�X�����q�E��t1���'�et�#���M�^J�8>���e�~\���\�=(}����Scirb�䱱�422h��3�����~����C��R���>+�D����~��	�F!C��(]��Zފ_0�2��9�������q �ή.ѝAGћ�pD)��"�_(��(0�ۣP~�6�r���+�����?�2PvU�.��������Q�Q�s�s�X��q|�,?�2%�Pn%��ryM7��`��
@^p�
z#�*��@6������_>K�7�J�����?q�	�$K�x��CIC�������Ռ(�>�����ş5l�C(�7�SV�ezT p���A��?�RƚV�M�[�d���9���ʋ�Q�o�ӓ�t����}�r��&��?L}�v����1+-,���9�&��%R���f)�LS#�O�� D���;�U�2�������M�}���__����q��@D���r�z�������t��-/K�I;3��"��hLͣͨ�i(4�E�ptvv�v8WĞ]�H�����v�ݧ���<O�|���u��@O�k֔'O�nJ�v~.=�?�ځ��J4?���	���x7}���᝼4�^婞>�a��ݣKJC�"�'A��N	�-�&��Q���;��=���_(X�3��#�x}?��D @kN�`�)�&
�z�⃃�Ӵ��'��(R��s7����wBXD#MEeG.�(Yu���u��^N��EO�KX��P�21�Eǡ���?��旸��H�?zӣ�?Q]A��WK^���X��� �?Ň0�c	KE�U�S=:�~��pt)�CL�E7�˳�:���?�*3������Xu�i���ߑ�V5}iL���:���U�Rd�7w��Ɩ��Fڒ g��Fn�z�44����g�Cg�Qt��K=`c�	�E(�p|�C�����H#\�A�7����դ�'[�(�*�ʸ�V|��E$��g�C��P��}f��і\G�KS�S���;j܇T>�ikg?�|���>�O��κs}���y$�ZhK�7!C����J�O@�\'���R���4V��b����YV�,+Vٖ_��^7u~�N
�!�Zf��h�gn��6P�Jǔ��m��׸e*��,��hI�Z~!���kzG)�E�b�4�D�|���C��|(��t�D+�שG8�i�R�Z,���DrS���;:P�;f�J�'r��x5�#���|x�4���+��^����,�W���,���6��7��f���ֲnQ�_��DFdG�hN����a&�y���!��<��0�}�N3y1�9/B�_%g� �1K�-�P�!^�=��N��l��م47���$��ґd���>>2���9ޕs����Ç��/�������[��R�@��x��@������>{���눔�16�ݼ�xX���e/^��l��-�A<6|P��G����N���P�0��T��u] _�QU��Cd�[m�WyPwPܡ��}T���̰�I����$pC��K?��,oW���G'�՚�����ۧ�����KQ[O��^�@�)w7�J���8@zE(k(��8��vz)��X�o�[E ��y���
�$��	5�)��nm��W�ޔ 3������=S�������P���vr���w�%�R{�zgCRj�I?������M�����[{�wɊ�wT7���>�~"�٠�h'��Pj��*3/�q7���AZXZMO��L�sKieU=")\�q�<���C@y�͒�~)5b�Pl���됰a$�0Q�`A��3"+%!H��2���=��Y�Q�Scӧ7�_�م���O���>y�~��/Ң���4�[���������!��
,(���T
�*��n�!����3����c��1V9h�̂a���Aq�v��F�d�a�0g�z�c����Qz�1ڄ����]�Pt�q�RȈ�lvÒ�y 72��^��ao�X����8~j[<�Z������ߨ����͈
G�p�LggK�PE�Lc�����eO];>�&�u�b�'��V3h�.GH!q�}�{'i{��k�����ᑾ�f��]��E|p�r+��\�[76f�� l�X6�)8�R���ǃ�r��)�<�<�D���Ԅ@S�ڬ
31����;���!�We� �n(��;�i��u+:�;kn����X[���@����=h��֙z������Ё�x��:-��	|� ����檇\a9[y��7��p�'���E+�2K����G��42��? Y�F��W�x�H|������v�_���.�6��j�+)�jt�$㩻���h(y�e-6g��әy(�0J_(� �F��k�e!���Dx�)�xـ@���(˯�7��o(<�w��#M��(c.�8xx����z��OyR�Ln��WYF��[�D���ɪ�d{$U�q�t&��g��7]�� H���&��F�x�ޡ܄rK�0 ��#�Nؑ��xy�J,�r/�R���s��z"ڹ�Q!���6+BY>:�M�� \	{���Ή6��ۓu��$r4W�����Q/�{���ts*fpY���Y*�S��|��nx_n�*��P�η��_+`�]�dz:Or{p�VW7�|�JO�H�?K�+jG$�T'|{�l�ڇÃ-��Y�No?�����4}���Vn����,� ���{[�i�eϞY1eDzj"��J��d_BVn��%�U���f^"O�kԝ"7z�i���[n���`;ܱ��٦�����*�(��#]Q��D�PnU�U�*�V����Q��3��D��=C��M+��8�r�����oc嶣eI�-#dD��I���s� =$���L�5:۳�������iPt�
B��ƒ�EcB�ȕ.g^u�ӭʣ����� �b������� ��Z����ӫ8:䋵F?*��!�r{z��k:���Q��ߓ���znC��ginf1�����ٙ�tp��z���[�Q)��L0e�B��;����y)jNB�M�&ܜ
z�m숩$�<�ӥ�M�E�0�����h�R��52�5�ج�A��ڔ"�^8
���?���S�UCB���m�Q�Q.C#�ibr2ݺ{����mf~;��f�o'��w�[��s�U��[ʍ��;b]!����Q�+#^��LlhA���S�(�NL儂����������5��*���8�P5&GJ�G�,��:�k����Ҕۃ���훓��b���lG/�B�%+�����7O����+Q���9N+Rhg^-�o�y�f^.��-��2-�`P�V�F4�|�b�Q��40ؕ�0-�R��)���-g�z*�K��A�B �+�����ƞ:_�I[Y����s՗u��U1��j��ʭ�?�� }~�o��B�O�o����s����,+�D+�]~��OYＯ�I�-�87�Vgg�*������y��e��uS���Q
�r4��]X(�	:���tcW�:��W�_�5l�8��̩��@�|RP����L���&c�}���^¥����7�׈�<!jr�:����w�Mqq��504���7�)h{:>mJ��gi��\��%+� �8A�G�*{��5ߔ΢���C�wP��#dt4�3Y�:Rwʁ'�k�!�^�y�Ju7����L����.��u�ķ�]��w~��64a�qF2�w(�N�N�������#ud�������#���N1�'+�J!� ��6�%�@G��"g}ځz%���ɦ��/
.��h�����>>f��mp�3��q�.(^���LO�j^��&�8�pq�{Ў�(�o3����m�x��i�	�#�!=����ﾕ~,]�έ���,����SЊ|����Ƽi����O9×����[:��7��Hk��=}:����I���>K/_̦�]�<;��`]0�0��K>������;��?�G?K~�N�yg�49q哑[)��RnW���vX�ܸ��ɛ�$3��}7�2rˆ2)������W�rtir֠�e��^�Wy+u�'�3�h+Z�V��FJ��>��%�Pϑ=Ж��V�ۑё411�e\@G�v Y����4m��,�j������w�%�T��H���#=!1e�*�@cz��(;:Z<:���]+����W�t����΁*�v�E�8Vo����اT�35��Ӵ�q�67Y ����L=� V.��a�T/ #!�E5x�&2zl(4L�OJq唄Ã�4�<~��g�Y��&�O��#zG=f��nvQp�9�Y=x�io��k>�\F���IP��7� �y3g�Х^2k;�$���Ȳ)l���R�z{���(���ʹ��eŚQC%�a�@/p{{'--,چQ�Ը*.ΟD~l����m�s=-�w��˨w�tyQ4w��p8�	���ԍ��iK|�#B��ҁo�L҅��������ٽ*zfb��~1q���{���ad$�<q,����:
݉��mU�Pz؜ŚU6�k���t��Mo����FB6�vw�~����3������`���ƺ*o&�7��@�CU��-Fmw�'�.h,��o*'�-��	�.km�B����45=���x�wo*MO�y� k�X�5���y�u[̈������d(��7ܠG�y������5��D�+�V�$<��r�K#PT?���+�Y�����������^�J���t�b���DD��)T��Ľ�UgO2�5���� ζ�[�T�x�"�W����2��`�����[��tH�uئ^c��t B�xַF�"����3���;�����k��)�R6z��7�S��-�����7+mz� ���'ݨv�c)G,s!+<��VZ-k$�Q��=�s���H���e�x1fsY� 'S�;O~�?������5㈕/H�N�)�c�.{#n�K�TO�&�զ���t73q�����c��hlH�/�%{h'9�[��6dPA~D�Dk�a*�����)��g����}�]irbH0�����,��9���1�a3�Z62K��3�ĩ?�!gj����h���eޠ1��������k����'�_e�o���7��n��'��2���F�[�&}�
'(�o�A9.%98�7�3��G�[�:Q��� ��qg9B��̝r@�`+[����ò8֪CF�хX��bˌ���h#2��;:ܳ�c�'��w���X�����R�E�1Ӷ��/�e��vc�-3��P���ޑb�`]��/�py.ev�@��]�z��� ��<��׈�!�G:�;�	Y���BNS�C���R;SO7���$gD��A��[�oєٝ����_>������׿�CZ\R����
%D=*�^3�<��㑀;=�ⷥ��\�k��~��_��4�]a_�\J33�R�V��v1r��ȼ"��tb���܀6���|Z[]M�{(r��R�� ��@e�� ����u���?�?I���������m)�_|�M��������c�y��=������/�;�=���2��+(�(�Tj�^)A###�U�E�ݽ�43��f�Ӝ�1jGg�)��F�^�
��V6�#E�e,h�95���R�eH�e�z}]����Fvt|<MLJ�u������E����R.�n�N��iT��3�ǲ�_�f.��O�C�"-,��mi�ܶx�ւT?Rz�0�/���8��v���L���^ZfhR%�Q������e�^K:SW7����Ⳉ��Eq�%��(%:��z��+R�U33���޶g�J�}���G?x/=|p;M��(9��N�;\���)R�Ӧ������T�M�4Ȼ{�iiqӽ�O?�:=~�*;ZQ��Q�8�F�2-�.*�+���]�r;y)����K�w?���}7N�� �_��).�d�� t/6i�C$�4e�$aqe?}����o��7��o^��T�:VC���S� bB�0
%ł�J�w��)��e��^i�0�����^���#iV#�Rd���NU��Ko�B��u��Kº�Iu�O��i5��V8�8�?H;��+�i}m�kn�*U9���D�y�����!�,G�2��A��ͬ��H��{��,`&%��ʏ<���т�Ey|��n�~ŭf���)u�a2m��%<���o�O�5�t��J}UD�e�3lhed�o�gK����U���Kǧ7���AZZޖ\��ޕ"��n���n�
Sxt}=E��X+m��\4^���Si<1��# �Z��1���2�!�(7�s����:���O&=�ͩ5�d�IN;�.'0s#���8�*�>\��<����XI/^-������*g3+}�Mf�K��o�8]�\m/�Q�[7��{���U/;��V�	PdY�y���xږ�LD�R�zC�u�V���˙�����U���cH�|n�s�#�|!�(?An�I5J [~D����!�R^��0Fm�vo�\c"l~�(E�!�\�p��������h��G���6a�*��v���7����:fp����'O��Vu@xѮ�IH�J�yD��@6�6�Dzұd�@���	�	���J_~�<��o���������S����Z�]�%�^�0>֟�{�GnY�0}k�.���B��Q`;�iU���/�$�α	u�nKo��;��M�˫�ի��`Y�6-���V��2�N�x��`�!�-�����(c��?��#~2/�?�gY-��w'�j������<r�L#��:3ݽ��:�j�N�ol����?��\[ߖr�� ���4� "ii�()4�l�:=�R�c3ƥ����C�Dd�rwo/={6'%�ez����"�����R6Ғ��eӦkr[YޒB�!�ʹ���)|���g�+��(�5�J�Ʊ0����f����woO��i)��"0�����b���βw.�j8����ijz�=,6��>e[L���6�����H�����!�^X#CϏ����FA��)�(q�#���moO�{���|�5�����^�#��u��ڑ��ԃR��&���aKi��Yʡ�q��-�6cKJ���N���PyҸ��S���J�pPٖ��hh�.o=���R�D"c��E!�h�-��#bZ����7%�o�Q��H`31�]��X�mv�2����A��~����Hhm�o6��Y�H���Q�%L�Q�61/#�ہ�#�펑J*�,���QRcsk۽ݽ����JPl�Ҭ����P��'G�;�NJ��,#�xUy�Fo^j���[���`�_��`s2��GR�Hk_��J�:l��2���¦>7�p9Q�?�<^\����}u.��<��`YBKk�
De���ab�c%�B6�Q���]�s�c��:�=���G�,�2��@5ad��!�KI����0=|��532�c�߀��Ҡ�h��"JQīذAA4 _w$P�w��Rg�H֢�!�wd�3h�B�
@�9��v����y���]���[>���Cq�U_��=�<����/�����
���ȸ��av��])wT_���Ą:���J-���iA��iO����c��Q�#�i��?��f0E�fFO\�I+F02�k�2��7�!�P���gdtHu�d��[�oz�#�!�Y�o�gwb�gx�W�u=�]�q�#��3@��,{�Q=_]]S}ݖ,b�1v��t�"%����0Y��urrX�������:�%;�%+�@�l�(�D22�g~ʨ�O�M�� O�O�	��ig��6={ʉ$���v�V����@5-V�g~�L���^:c'�6�\P�nr��.�~�?+�tp%?����w'=�,dy߫W���yt�M���{�ʆYc���r))��,W����A��e�����XJ�M��rℝN�Eu�Y�]� �\a-\���@�NP߼�T�yk[��^�G���c�Vz�� r��]��od�u�>Fw;�Kw`��u�e��h�3 ]n����ֆ�x)a.ס�1l�0�>j�Bʁ�N��z��F�G��q�I��! �s��X��ȭ�ɯ�))�����������Y��/~�.eeh��R�Pf>#O)
$�OO�����&�j�܎�Gx��)a
�Q���z.x⵮�[�VZ7�wҦ�ʳ���
������zZWv[����MH��,�B��P!�7���Y�q&)g�6K�@�X��Wh��	���="��ɳ�!���q)?���S���7���|�JxmX�B�q��&��c���V��Ԍe�ƒ�3>�K%JG���S>RDtb�1��1b���	J�QHL�1�4,喍�L�_�2�����!�I5�VnE��m)�Rn6]�X� �x��
�<�MY._R��У���-�+τQ|3n<Go�>���W�ybQ����*_��~�)�{k�Pڈ��Ӄ��P�ͥ�n(����E5�'j1B>aϱi�g�e�2�w"k*�$��ᖥ�������Q�S�k!��p��x(�yE�ݔ�ڗ�g�a��)OP�ECI�Yw�3��pֱ��	��z
s��:�����B����ι��������t��p������W���Q\��Q�-n�5կ��^��ŕ���+�N��Jɠ�c$��P�T�=�J�}�P�Q�ؗ��0!���oA�	+�*S�_�c����A��_D��p�;Rn�ܙN#R�X2ҫ:�!~j8��sn� �C�Rjc��gp�3��H�,���H�L��0l�dĶRne�?���ȅ~���y����+�|�
�O��s���Oכ�G���s�b#?q�ED�Qz��ɡ�t������[����Ko?�L�;ey��ٝ�DznG����:Nf4�9��	1�W�b�D�!>�b��1Z�)S<��ݨ�����}����l�Ga�U��,y���" �Ȉ�YJU�<�-d���ی����>�餱T�G�#�O�d��F�R�6�\�@���l$et&�h��7�Ss�q;;T�� ���Cu0X֤�r_�lZ-�������b��Q������Ȏ5�G{� �� ���]S�	?��+����7 �UN���U�ǿR��������.GQ7V��� ��3��������S^:�ƹ�������433�D�e�h�H��,wGd�O���F���%�&4�OE}Px9�k��L�TC�����`��Yi��mY^R�Fzt�-&^/��R�F8�o��[��oJ_VǱKqƦDSC��*���v�8򓥌Qf,�D�e)#
�j���WA�r�J>��	2;�6a2H�i��R��]�6wh�?|�� /J7҆���?�e�1�,� |�h_NL �g���f�=�I$gGl<Ѹ��bZ�(�@1�nŕl42����������-fڒ�-�r+�{cU���U6C��+�j��Ӯ
���8��d1 �J�� ��F$6=�X�PŠ�Z@��9#��B@/���G� C�e�p_�BR�!c�Ԡz�ݽ��%	*��9��5=��^���P@�U8��M����u9�J�r���L�X�AV�/i U��J�P���6�f��U�
� &�N�/�%�rg��ʫ���E~-�ԽCg�@�EO����w*�GDQ8�6��.���b�<��8==V�d��+	�R2�T�wSG+ǥp�q������cv�KA�p����^ۖ�&��5׬S:�2� D8�d��P,��l&={�<�|�";�IKsi]
���J��\OG����h75_��i:N-��/dؾq�������*�*Z:2�sF�c���:<�,�_�2�������l��R=��eZ��U��P�=	[��9���ښ�y��QXG^bA�'"J�|�r�zmr@�(��3B�4ޯ3���{%��M�Oҋgo��3r%:p�1(�����,=a�yA�Tv����`��c�ǉ!���X����gQ�U9=*	��%G�_��,E ���Q+\"Z�S<��Ư2�0u՟/�F,�!�ꀉ�(�7},�F��w���,Bx�
<X�L�JV`DK�{�ʠ�k����Ԅ:�l��Qe�����=ӦN<�T,�]����R����H���!��F����o����j���i3saŔ�?�/����1F�8N��v��o>�0:����3���03{��`ooW��Ǳ���dV�b��F
kK34g��P�g8Q�P�mK�Ź��Y�߅�-�i,'���]��G��{�k�O|l�U��>��>�W�dnoW���˦+�W=�`�E4b����g��KF�I�@F��}�#9�#<��?�>��a
-�U��zU^$&�Ku��E�U�]�&�Gd�x���2�v�`��d�3ۧ6G���.�@m	J<a��e>�̠�8:)�ؾ:]	m���ww��,�I�mCƁJ(��d�p�f?�@[���䔏)T!Ӿ{9�h�o�L?��!�
�Tu�g@!2����)C6Q�ʻ��i|��9�� z�����[y@��<(� �R/\+��J�2�^�|9o�2*F�8�Sl��,Z���CA��AT7N�X���XIb�:�QgV�q�ѹѮ��u���[�n�0���
`��)�)\���9F�˕��K \�������~�����!ȬN2n���Ŷ�oЧIh��7���%�i��z�Rn{$Ȼ�kBs��3*(S�bn�ѤJ�;�%�8���$��T���)|s��^)����`·��ie�>@a`��I������=jԥ�w
���p�]�$ԂN����v�/-? j8�NUO�b{�)g�z� F���M��;�@#��VJ��,3�l٣����^�z����k��^\��(,���&#�_|�u����ߦ����N��<��Qn(�����p,΅�f�$�O��G����V9cǣ-\"��(�Y:�?V�kSʬ�5{j$���fx��#)�jH��{]-�m�����x�q�Z��ٮ��o����S|[����%�z_���L�♔�x�k��0����4:<��''��Ą��%)�s��n0��� �!�*:�,1
F�z`�P�ᛚd�̨�Q��\����`�ҳ�:�w�!�!��+��܇Q�E��V�t�ٹd©d;�9�H� �+(
�ej�;���ru���ˆ�J��;Ȋ�8�#fN�?T|Oo�ܚ:-��k>�SXC�,b�B�Pe��D�M ��T�W�d�A��u��w�^�>��~Կ
(�R���J�@��OHY�Myy��V�h�����ю:R��>HO�>bJ?deGL1�����	cD�ҡ'g�J\tp�Mgeԗ#�x�����+n����ˊx�����
7~������iS�"	�	-;;���̒�Ռd�B��_�;fL%3�%ǰ7���jz�������S�mgVh)m�c��}byR_/'2�h�����Yn�2���֝�	?��E@�� �gB�xey9--.�ٹ�43�B�R8��l�yiq>��3��#x�*oH���T�7I"�@�)JYʌ#����X�#�q�'�j37��I�g�*��l�q��Z�7T�%�<˪��6��~���l`�R�j���/�"{�C(�ʃ2���G�+��O�)? �*u�ƙ��n��?�
�dE���G������s���&�vu+�8n�{[���ꆼɰ�"�s�*l��`���� L���3��ҵ��z���O� Y�(���S�2�r�1hU���f�4/CC>���SE�*o����&�l��QϩWЏs�O�, [r'2�Ce�4'@�;�7�.�4�3%V�=����!� D�q"B��st�$b 1�oGB�8O�e�ʨ+�v��!%���g�7=	�������(ng9�J�d:��[����d��x�l~`=�����F��72 ��1M��)T��8�F@1��$�'���z����DOɢK���g��.��t�f4P��Œ�����,�`Z�GU@:��8�#��b 1�XS<�^�w{���2U�ȗ��l���`&���(��[ieE�yi!��I(ʭ,�g��<_�x�������'��o���ͥ=);`�4�=��wW:�T�H��ߢ�����!*���r�[�����U�kә�Z�ZS�z���i&�w1�'E�Smޠ����41ғ&��i\0*����4��!��#�v�A=wu��lmT��8ň?Az;�%����GAgz�S�̩���
�����6����/��v�t݋�=��(D�!L	�?�5�}�У�+8�P ���� d�h��k��3|��J��J)b�k���{��I���o�_|�����R"�C[V��[���6�/g��(�'�Sǌڊv��
�:��}[w(i����l�Oz0PmLˆ�MN�5U0⪽��o�����Px���TY �*94�;�{�����M�_<OO�?OϞ�H/T>�����e�&2��&��C����D[C�(�mO��0��W)킢�{�C��Ώ���Pp]P���j�fw�
釼�̕����}P�1#y��#�^r\��yɯ5���k��<���L��mI�]M��KR0�x
����=ё)讎�ԧι�au0{����a�)� G�1���:�/��fV�%(���e1-H���}e�����4??kٺ�S�����a�ւ#� EhB��t[$��a	�������t�֘�ao~�f��4${d�7�p�����Ҩ`d4�%w������$V���˃�?�8p��s��W����G�	Q9sr���g�!oBҟ�ʬ{0%���ݴ��4�����4e�-��t�-���!3�˨�G����SV��WB�A!���l����@�h���_�Ѩ'ʯ2�B|�΀1J�@ i�4�7������s��:|R�;�\�r^\N� �T��ej���G�s�7X!h�#'!����GHaH����z����ŔJj|�[(�@yt�^�b�҃�FEe{�2�n�כ�)�V����8�QS�	܋�7�z�F��Q_BM�"��o�f:s�v���l#RpPL�Z�)̑�Ψ$�6�.��$>��HU���i�Ǌ���K	����Y@�ܠg�-L �.(��0>�e�zs]0��P��x��$�	�(��HP3v���}L0�L$n�y�N�V*7	�v��te*�)��=�L�p��AX���#'�#Ew]dye%-�ϧ��)9����R��=�r8���!�CX�<���)�,�PjYs�����}�H)J#Cl�O7'&ӝ��ӉC�ـ���)e�������靇�ӻ�ny�ɣ���o�Io?���~x7=|�n�{W���w�=��E|�-~J��o��S�R^{�c�W/�x��ʛu׽=\C[6��(?tL�#T����z��*% �p>(��^}��0�$/�Ѐ������w׀BT1:-� eǊ-�|q�JG�揙����>��_�U��������������������*}��/
U�
�#����u�4}@��8Vg�H�Ng�MOp3���!�w�r@t��s~%��?� �y(��a_�a����\=�DbC�qF����?O��_����N�������7z�m���/����d�-2+��q�z�ĉL'-�ߣ`�HQvJò/+�up;%�6Bʊl��(�m����j�w���sV��|׳yX�����!?�b������\z���/bC���e�n2�L���Qe]�:a<on�q{[y�4����ڤos�Q��ݥNs3t�Vf�y��@ϜL���$X��3L�_���������|�����Ϥ�Rl=j��&�M���S�������3!(c.d�	(u�Dp�M)e߃ l�}Kr�'?�A�ş����~�>������?�����ӟ|�~"��c=��Gr����L���~�yN�`�Q(�*+��1�5��k�˕v�m8��ė�pm��ye՛����,,̫��Q�'��H��9�h9����e����ܳ/�^�'��se6�w�1�!��2�	xV8
+
�ҿ�e�?���~���N�؍_��١p�d�<(�^�^l����I��� <���w�E���ԥ���@ �#��Z��y�De���@%��3a�!2�A?C��c
����O'�/���R�)HFC��P�x�MQ�7�[&�(X#�H�8�(V|c�
C�L6��G�b�0�G!L�R�NiΑ���p$3���Ʊ5m&���$��0r�E�"�$8~�K?U+�L��8�/(����ic��=�8��������Nx� XDe��?��"��69��@+Y����x<��Uv�i?ʮnu8�0Ja�nfS�ԑ�H�c-2���M�&�d�b���3��T��<	������NW��,�hPN�_t���#�#eW��G����8���c�n���z;=�����w8�aB����)�7S7���$�G|��;U*?6E���72<������B:-ތ2��rg])�"��\��aTɼ���|/\��>�r ��2��	i÷댢��6%�l�:�ѐi]dF	lY	��+�k�:Mݎ�(�p#�4Ϟ=OϞ�Hϟ�L�jX�]]]U�e4Ԗg9z��+(ߔ_�PiÇ���q�|Ic����)!�8���������r�|s�G2�3R�h�Ը���ɓ'髯�J_J�e$����� ����8m�2(3�4nV��7���Mм�z�L��N����P,��x�u��1��WA��%��Rn�I��rJkl0E�a##"���8��S홤S��p���!�9�-#��/\�~�Zs���wFs��ZS_w�����V��K�mj�EO���+�K'R\+��!�R|�8;���֠&x��2ϰ��Q�^9}B�gf�j�%��sA�l��G��������>��駂}�����(���]_�������)Y�	Fq�MLW3J!z�?��x��D����Q�,���rf>�lyfV$K�'l��XЃ�}�h��m)��Țk6��(�(�>�P|�Ag�d+��-Y���Y�>�Ii7�l�[)�6�|�f��ʪ��]�)����@z�z��f�(�QÔ|Z�s��">�E�!r'Bگ�H[��n�9m�cг�4"�'�&���#�D�h�����)�g��BaU��T*t�bd��;X��k0EA���w�"�T)��Q���1H�����1G&1�HAֱ9�Td2����<��<���5��^�
��X�3��ʥ&��*��4��A��t�o�#N�L��YV�`tP�j����η;uHP���!p���m��rHU���pc� *�	@���F�q��c�E��hX�n�����y'/9P��h=wa߾{+=z�Q���~�h>��8m����{�?�Y������������r���T����C���R9r���%Ӝh���`�3�	Ⱥ�����#��Xp��V��n~��ӗM�} ���魷�;�o����4:!ExrD���3��F�t��0����谔��a�@@
-��Xn�Џ+�������rt
{�������[YҔ���ƀ���.)�aQl�ӯ'  ��IDAT�ӥ�¯�,�(��#���(��� �����u�x�,P0ٽ��B�#�QL�>�*͢Ѓ�ؤC=g��!�͞��'J��)��!�K��S�ʻ�G(�E�u#-\�!d��o"��nm��u��C��<� рgd%���n�[���H�p�����yt�ʤ���Ư�B�z�Ƚ(���e�\2�^�c�g�L��(�n;�~(��+���VX��Em��+nr�;499N{;j6=U�LbG{�O+����v)�¡	y�PX9m���ܞ��T\��iͬc=g}�:ԭiP���@o��q�EI� @�c�cֈS h=X�t*�u�>6Orsll���cF�i(Gʁ���n��Q��_�ssU/*x���f g�2c���T��ݻR`ߖ��A�ُ?L?����c)���(}��#�o�|�P~���[
sۧ+u�~�hQ���:�Wꕁ��^�̛@�\��|
��tv����~S�2:��R\�f��Q/�N< s �
]c{g�{ 8E�cP���N3�$�*��C�y�^�}>U�<��ҭ\q��o�S�@��6P�X��됫`�Lpl\%%zFg7�9��#~�_��%�qy�i��G�;!4By$0	`�,E�@  � xH��cVVֽ�hV���h
�&�/N2P�$H�x҃GYl����71�Y�2FzP�x��[ ���#�X�'č5S4�;RV9
��Y#%��QVp� 	a�^��]��0��B�Rq�A"�vVd���	�YQ��\�@�+�U�Jߪ�È��F!ɕ��0h���&��E��^&���lgFOٟ�� �����;^.y�ᡌ/��i��Gʨ�R�5�[N����|�i	����.�%��	��޽�>��ӏ~���λ數�i���c������=�e0:(4fB�x�@YPI�t��B�5Ӯ��)1��]b�#挪��85B\�<:>d�OWG�:r��"�R�:�|�3�m��q&jxPjY�4&��Ux�A�(�Q��{��m��E�ş�4/�˂z-�e2�R�Q�D�r�X�s�	��2W߯3%�� �OFW���2r�l�O5������xCCC���I�>L�=L���M��P߻ܘ�Wo2FOyǏG����A+���9�X7�7 ��e��4�3M�h��x�S��/Y)�Q����{$���|q��D�u���8�fWY�I.(RA��U����2pQ��S��H��z&��G�c��\v�Aq�\e|j�J'��ƋW!6�^�Q�3[|-{<�D;C�Z�N0�a٘ʉe#��y	R_OWe�sh����t�OS��0��Qw�C���Sc���d�}s*ݚ�|���,[r�TxЊ��sj�ݐeKQ,[�m���G[��-u���F�l����N�Rʎ͔Bϕ���b")�(���+}�%�!�\=��i\��,�I)�C�2
L�1�������w𯃃���u�c�nʛ ����[T�վ�^̐�T��89��@����X'��e�w"f��#F9s�V�� ;�����U��W��l+#���A�o�bJ�~�A~(^��q2�yv����K�r�Q���\D^�d���6�+��2�2_�'�+�@�q­�1��f���	?�� DC 7*a r�IPI��������{��7��z��qZ\����aŕ��˒Jt(�b6�۪�$��OvQ�`b4vԡ��C��d��dPv&��&�gF`XC�g9�R�p�)%�װyyM�L3(og���!7���be�v��/;��"ޅ��_�am��l=*�� ~�RBI�" �G�� �������;�/t&�T<ʫ,K�.�y�L���\]�.�����b %?�Rٯ5��}��g��Zg:"���<犝���pG:��Y	{n5Z^�6p�K4�'F��ｓ~�����o��FǦDϖ�����=�OϞ�މݹ���V	�.�KN�a"��#u�v�Z��b+�l����S0_	q�Iw�ʈ�;��jhԑ���J�kiM���l�aڋ��l���A᤾yy�%�y�>����m7����&\��FB�	ᑩ]�N��W�FM �R.�绌�$��5"�ca����s��4�/�� _8}=���ș&74(R���>��g���៧_����O����;��Q.;Qǁ�u�q-ʈ��, : 2A����|/2��Ӏy+�������IÃ�'9)�2���[�W�H6>1���v���~�����?���I�g�쟥�O�i�G�����{�e��d��/T���u؎-���D�pe��e�* �(;�a\WD�SFۥh�3�0/9E���u�up��`)G�:�m�2�?<�k�����2�N�s6��KJӐS�`����Zz�6��1K�Q\ix�OJ�p�-e�����]���%>�"	.��R��
ޜ�ɩ1����5�����m�~���D3��:W��Y#�)$GG���й���)a!���g��'O�7_?Nϟ�Lkܴ�8Ժ*�iwk7ͽZL_|�E�����o��.0��N�^�Z�y�+:��el,KՠƵ��A�P���&�V��h���P�O���ٱ�c�v�4sGmR�>�N���t����Դ;��?���܁����tG$��p����cw��K�SY/n:�E� ��N9Տ��Pv�=�/��e@��� |����o~��ϖ㼓�P�j�#��=S@�2�k8�����z��
������j�<ؓ�ឮ+o��@��4v�J�:����ͦ%)��+�`oK��@�y.�=�{�9oW�{�I�Kwx�P�l�RBA�>
E�F��K ��@4�GFC�E���?����PHa�����,$?9���������a�f�?K{{�ikg_ʊ�6Ty7���֮�^)S�R�PFO�6��*~��=�2�r|x$�70��W4��}�����9J{�6G�鈥�_�urT �I&
�/��ܣ��gE�
��
�؅��b:"{����)v��(�`��l0�Rr9��[��J��F0���w�$�x1����i�R��1�l�"%7%��E���������:T/ҋg3i�v�kp�#� �Q�jj��/hAg��t��hj,��<%�Q�T�ҡpz#����Z2�O��ơ=	�C5�'(?�S�Y�F�xQ��!�#�̵�	�(?h�dmS��_pR�`���D���k�)&��_�s�=�)2\^������E�1T&C�M�7ӘgpF�ⶾq5:4����I����������z��D���#G�r�gy�G�����f�!l�P�����vS��\�Û�?��ȕh2��Qɢ8g�G��h�����G���x��G���{n�9b�8x-�Eae3%~ܱK�1Т��q�q1��� �s�������� eR��e����n񏺡__�W�Ƚ�	�섯�G�]�o/��I�@ݗ@���['�3l:S'A��vu���?-J�u��RPYz024h{��Gn�i@6k�Y�:�o�,[����*>:#,W��L�C/o��n�/���י�!���:"���۬�^[c`h��Xk��Q�����@gg�җ�K���'��_��Ws� +��1�sd#�N�"��W��@<��ܕ�R��� r���IyU�%O�u$4�-�]�^�ŅM��=*~g?��@�/�r0��ɩ)���w�}F��� f��_H|�<�ݬo1(�M=�Mߢ�G�+2%x9���?�^�H��-�Rm��.�ht&� o�n�ke�&����VR�/~0%� ��+�����Uyq��{�3-�C�� �E#d��?VF�b�I����`14�aN��S�"k���v���Φ�yS{[�8�z?�r��ޏ�6U�wD`�䤫u���!o̙�T�����)`*��b�,�/�y�zP�&<U6J�dԾ�l�9�G
���O�͍Q�]-�$ĴZOp�G[}���nZY�J��G��/��Սm)2'VHw���ڑ�H�ݖ��}�vv�X)�;��w�oKJ��^Z������H��[is�c��IJgR���!%M��5���p�k��x(7�W���e�j�	��H��7�S����,�+�WV�-�P�sЏ��(������'<��	�_�{ KKʆ9�.m��]g^I~�~��ߤ�o�.���+ٿI��>O������_�o��I_�,}!����&��y���������:	�#��N9:�����y-��TOObD�F��S�C�,W�i&��p	�'o���#u���쩣C��Z)���N
#U <�����C{����w����eN^�zF�f����|�Q6j�,����)7�����R��Nع�x��<3�,���AW��,��{�/ �+����N�p��M�R4��+w�j-1���WN�P�n����,���|��c.g�q/�Z�"���z�cZ5�����SL��z ���?y�����:>WM����e�NJ<�������ӱ��u�R�$C�I������TV���L�g	��F�^L���.ʬ����ɏ��.#ꆙ�ոR���:��tB�)�|�2��2'dgt"��A>"' Ub9�l�}�\P�� ��ܩ7T+M�9��6p(7I� ߉�Lq�y����)(#��i����6*���±�Qρ�>O��$R7`��:���LYO�)�0u>�'D ��Ln�dc�G���Tf��wv|"��f��O���Ɔ�ٙ��d��Rn�������K���Z2J�fn�cŌmi���+x�g�:��(C?2Yi7�V��U.�����������=�mެH�������Y����Y�?<2�%
̠1+A��?�|f~���R�I{�v�Y�(���M]��E�8�-䒿�MP�*���/��wˮFD2�0�&l�q�!����߼)_�=ځ�e��W�qڢ]�X��$�9ʯ�]��fʌ@̨D�y�^;o�N�5ҿ΀{��!k���q����X!�P��a|!��E���XKĎr���= ��	GU`� �~��Yy��O��߾睔o�}?MMOx�7xAO�P�$�J�a� QT��I������7��L@,n�9��:9�9�1^{;S�"�t��yRB�7���rz�r>=>�^Ȟ��r��ʫ��b4��-*������meu;-,�+�rz5��^�p&��W��r�ք�T��yGV�% ؝W�zw�+��E'�d�d���*74BxˏA�W����S.z:�l0򈐕�b�Z8.Ʀ£����(��=ь���������͗O�g�*��W��������gOҳ'�Ҝ:+Rd׹���w�{��#�!��������R�9�����:e����I&��$���r��02o���b��`���<evF��L�ޮ��@S~��o'z@X��,�@�I�lt.-(��֬+>Vz���F��h����g�W�*�Vx��E��j�H;�}�.��W_�_O�*`�د��2E���N%@�!bC��/-.�E�
��Ae#�-8�v�s&�a7#u�4B]gy�
W��7�n�#v����(�~��-h�� >e$��Ǚi�$�Ϯ|��i�p&4�AtZBY~(�W�#:F(?{�#��؊Bi�
(@6��K;�7��L����7��w���,�:r�'���2�����T��Fĥ8�lΣ�G�-����p#�E�8�����ޞ���Q�#m u�:A�k�C9t�T�O�,`"�Ac��D=˲8�t \�oE{}���L
K����m�[Ir�A�R�>U@|��;4s�e`������F���^��+�*Ԍ�@�iU���d�42��^%|ؼ:��`,���3t��]f
H�A:~(��!�U��cO�� �C��:�G�Yg���(3�^.�K��{����d����2�+�Ə����ݰ�Cq+��|���V�C���O�=�1�5�.?��a+���r2��x�++�EAr�����:�����NeS$�hFǘ����u?��6�*�>�Jo=�'�v�{�`:ݻ����~�>G�|�~���?��O��?�azWn������w�
B�0����`[
�|�����o�p᭭=)I�
>��Q%I���>L�˛iff)=}6��y�"}�͋�����[Fs��Pl7�hm����X�����7>���/�W_?K_~�Lq>O�_��>o��cFhϽla[����NZZYO�j���ܨ�ؑ��fz=��Q�]�Vr$��LaJQ���&)�`�kM�Er��5�	n��z`�!QF"86���ݣl�`6�/�W��K)����S)��O�}�GhQfQ��&�����U�0�� �<rC�L��c���k�cC� �@�=1΅۹��S	�ݵb��Δ���,��!KM��DcÒv)w��Ti���aٕ�FFn�ܬ�*>:m>����A������K�����-�S�tr�c��ީ+��+��1ⲑը;���|�A/n�9�p�{���h,��<�ӥ[��7F���r*9Î��ť���'�2�V|���7�<V�����LC�m�r��+0��v5/�p���߫�����}��� ���I�4�|W������ŅEƹÿ��oӧ�~������X����9��Yu>���\�q���X��U����M�N���҉�.����ed�,���a�E��Eqjо^���P��~�L�:���k��W�/6U�6N�a����V9����BJf��y�y��ȤX>���,-��n�2H�e���>V�vz�B�2T_�-�_�Ђ<�֓HC�V0�+�"s�
~��%���l�d�ihh$MMӖ�O���I�����76?+�]�\�0�n��XĻ��GF�d��3m�@(��x�m��D �+����2÷��W�'�#=�[:��f�#ߐ�2(�x��BY����a����c��9ڎ+�5u��\��w�/��y9����V:֤��+
�Gg���:r��2\ ��z
�*�0�P�E9�>�����Y�B�z9�+�� �u�����"�����8�s�U�������񋯣Gxbd߯5��#T#��M/�F�]��955�о�����?|?}�累~�^����.���I�����+=x@��J7o�:�.Ur����ʕA�se4�'��P�|�Q �/�!�?�a���!�i�k;�=[H3�VԀr6wNo�޲r���W��ҋ�\����tţ��ۜ��u��R`��t\��̍5�譬,�.+�Y7��0?{�J�¢�^�¼�%
�(�+�ū���)��S)՘?�߹���&�c�䊤���$���h9��m� 0]
_�s1���e�MiQEQ`@�' NN)�"ӈЇe�#�Ci|l��'�Q���T�igK��谴�,���^sww�xmT�6��޹��&�g����%�D#�^�\@���㲻s���gt��9��3��P���;RH����d_
��IJ�gC��u5�*�cIƌ��5x�p�����Z��t_;��m<:f���,��8�������2�r�#�9���K����� �W�����g�B��2�?r�y��ͷ{pջΔ��k��yG8xZ|�N^(�-u�����W_}���ux~�i��/Uw���,��;V6�o~�v��hh���iۛҬ�F�+�A���U�����M!�j��!���(:O��:۪+�����So���~�~%���#E�w�O�H/^���\�|�KF���k'�ϙ%Lء�zTy�������z�
Sv�j<�x����S���Iv�}?_������²�uxcv'hm?�����g�J~��M/�]�r�-����*���k�At�u��d9 3x�Vr�ܒw:�J��?t������D��`�S@Y��4�	���4!�f+�c��};MݜN�㣩[�8�N!�����>}�J��Q��ᇲ�N���C�8����ݷ�l ����A�1"�_�rd�W64�M�,`��Y�qf6���#���dOe�R̹�[jſ+++6�����np���u����&�(�fiB��\h���r)d?K��)�;��"��T��4�y%��Dve�0�@���.�L��k�|�UC���M��e#�Z(�.uѸ_E�&05�Ʊ`�Q��Un�o�mH�(��6��G��3��?�_���d�U"w�������
H���x�bf�����4�U{��i`�5)�il|B����p�%���[7'�����1v}w��[�g{�أ�k����u$�P�����N|4^��W=!1�9J����st

��؀�μ��铗iqaILWv��]	�u)NR�^J��J�Y5�kk걉&Ѕ�('LC��b���:Ī����6R�P�QEB`�$�3E}.\8�l?�olY�ސ��:�;G���F�����������Ӝ[�����A/��BKi��=IK��iiy+-̯H���$�$h}V*�	��ʳ:�F(h�W@o.�\�����)#p(��1K�MI	���1�&tg5����nJI�v����4��H@0��i��<6QP�w�L�St3ݼ9��{���;;({��!Z�����ذeNc�T�C)�+�{�ʹ��bA32ܗ���RgW-S:!7�Kp�v6r���k�u`c�񝟷��N�6�;�)c�;%�Ʌb*S|sp��U{t�8��c}z��s�6�׮�:LNN�.	��6��Ql��miyA|��z��3�����M
ȅ����W>�ow{�`W�+m�7;ʆ2���[�n��`��ƿ�'A�{��^p��1W��(��n��i	&�g��"1�-E�@�%����V}��yojaC���p�`K��ň�Ϋ$aPڕp���w	J ������S솠�����U7�FB~�~oS�����_+<�
�ZcK[�3���>�rݷ8!��}53��?K��Q�M;����C��%:���0�R�2霒e�Q��AN|�
~�J2a\�~;dLVֈ�H�x,wBI&N8�����7n�<�}���H�ګqɑA�nlQ�=I+�kR�_����}rz,����4<< ?MRF�%�X���3���_J��ȐG:�cIK���=+���R��.���3xA�p$���lV:���#��NbQ������I���2�KF�vw=��t�׏��{O	��7P�K�cy�%���m{v�K�V��~����Kw��Iޑ=��FPl[$󚄋�s5�m>��`Xt�N�%��'���@ЫW�����4;���d��f透o���o�P<�q�\]�=l�i:s0�룻�����444&�.��$�u'͈_�������9�����?o�;Rr9Y�#���(�(��	�h��d�� oqN�����^3�rQ����v!t���5�[�#Д�Ԣ��t�����V�4�����a�}lx'L �-*�m�M��e�GgW�:�*g�TjP���C�q݈�6�T��7�y�O�8xݔx��+u*���������V:�)����9��(G�Ћ5��i:~������NS(߀0���Gq}&*���CXJ5flzi� ���Xpݧy`��G��� �6"���m�͑*/Gn1M�;~�R5đ�����l7L�{����F@��=Y !7?~�$���H���K���<������L'��pW���n��2"�B�t�1�X2}	N_��㢋}�s��2kwY��F46��[�x9#ܞ�Ͽ�2}��g���駟�o?��=ыJ�d��ʰޣ�_}�"[ Rl���i<es���d�|������ݣ���P(3����Ǉ��|V⣷n���>����λ�Ըܔ��S9��2-'g���[�FӃS�,��O���2�/G���P���L�����Q3b$����=ֺ�f����NZV-��Xr���p�,/$��T���ꈬ�Qa���%(w��a�/�6�$����]S���4��J��X$v�+��
kŹXd׍+B)Fg��h�" _J�E�+wF�<�e@(�Iuˤ
���s�c�ۛ��4Sޯ�����H���+�>�V���^� ��vE�C�����a
���r�)ߡw���_6`�]:j �����1��(W��PB���d�� ٤�
]�������9��	zb��F�&]�m4p��FC�J�ſ@���������62��0G�ѮP�I�=o��y�me@�\������?h�t>�㌂4;��^��U�a��Ԗ������hU��:t��[�D /ȗh i�c�/���9���R��SI�����jz7�?v��'��{�$����^���ŵ�rf)��]�(X�~&8���m)��R�z����Z�r;���=��*^�@�_F	�n^�7}v	[xz�J�a�
����~Z\ڑ����f����I�h
��-FnYj�U�t8X������h6�Y��f8�Xg�q��(���)/���l(�e/k��_R����+�m�EfY�T�Ap�(H`6Ԩ�@4ϸӶG��W��\�� �v^�?�W@1�R���⡐T�!4��	��:4����e?��?��Z^�G�~�@LLy:� 9�ڳ�� b�*�z�9n�޹l�R�98O�j�7�<�&uu�`'-��W��3\X�L����Fz�|-=~�"�rM��N�r��4�!�ѣ�@o�"`!O�!H�;�Uٸ��Ŋ���\��/�o�)�����M������!J?
��������6�O�f��#�RX�C���l+P���J��,#��
�i�J��#��p��ܜ��<=~�$}��7��Ϟ	�yO�Гwad�G?�NB�@V^%�b�3[�b+� �3�S��M&�U�R�h��X}pT��L�1�M�ix����H�}mijj0���[飏�O��(M�S�󴹱��f%��>���F�P/��y�%��Q��w ���eD�;'kOl������8�2J����)�7�(})��imc+-,�#��.���Գfn��])��^O��B�|#-,p,���-)���SĨ<4���2>������u�6%87Թ�ظs�dgWj��I�	ف�}���t�zzp��XN$��8�;�'|�cGLg5�{����K|'����	R3zq��g� a��������!����PÕ�M�#�5��V��G������_����?��:A�{���<�5o4�*^~��)�0�7�� s����h�=�n�#����T�:ԍ�!+~^(>����\�P�7'z1r299����u��_�������S�}�jX�h�X��N�ДR���.DA1(kFi����\F�����G��Bnxi�ps��_C�9q�`nO(�a���y@�pI�80��"���8����qآ�*M�UIU��N������M7�eKR~?y�>�����O�7O�{����if.6� r�'�g@�ܶ�H��]�t��(�\��Z�X{*�@]�(}�V�Cd�Yy�t�tBvZ�-�?1�^���?�~��/����'�7����G����Ag�Qę.��ǳ��O���~��_�.��(G*:�!�%;�W�:�����E���#�>>/^)���h���!��[9ϳL�A>f�Ї܁3U��P��H(`�N�^�6\mDlL��=�����+֧�H��y��ʞ�]�*k��_�;~�+�5�B�o�I<#���ܐ��A���M��Jl(t�.C�����&���3*g�$�R�@�A�m~1e���G��K�J��c��������@~����#_r�G��6��U�DNeg�
�襴�ЛTю�������rn==}�(�u&}��E���g鋯�_�ϿR%��e���U���W�of�k]p��>�V�1"�0�Ko�ę�!�Ja(d*�Sf�5���S�'������ڡJ�,�u&�uv(��DB�i���M��}RD����{w���"CAE��K�#>P���slW�놅J�1��Ia�/x
��8����#uvw&.5@��b��ЎU���F~�j���h�dfr�bу��?@_�d���c�(�E'_{��L��
ր(�k6���S(��C��;.Yمq�`����3MN��n�w�{+���n�ҙ��g��i�N������>���=:��d�,����b���f��F�Xnr.��?�^e  w����`7�)]�4��j,��G�5���2��N��2;�Y�-�wU���\x��%qU_�;�RO��A��!��� ���dI<v�=����Î��pXݢS��%�{��O=,�U|�B�2W�"�cC9�bpnE �'<\� \.�vհ�H���Ha����f���"��0U��/���ﲍ�~�D��g����o��>��_��:?o���Y9���+��������US��� �L�o��� ����+8���}�waFI�*�F��J�gLԐ�����(�C�<��?�q��㟦�����q��ޒ���Ҩס��	C����x7H��!�rل3��F�dEW<r~G����\L��uc:H68~�r�g��\��ɊF�z�e������b��e��'�S*���9�PJ���Vuʚ8zRlg�$�KV�I �O�D�ޟ�/��QX�b��lZ�3E���5��IJ����Yz ���r�D^��ٟ,CrP�;�6��e6T��4����Y����'�/���2��Y�(��\fӷ�.ʍ�+���]���NL)�O�y�r�PVW����'_lL>������Rn��~-]���,gB�@���t�hwi��U����(�Hz�	�l[F�i3�P4���<mHZ�[I/�ͥg҃f��,/�'�6Z�Vx��g����(y�l�K�ǌk��رǀ���/c�H��v�f��j�NGuE~�� IN;C���݈�q�'�і㖱0�Z�<����s���j�݀y�������<����/~ɑU(��F@�S�ݰ$�~�y��jW���wJ���:��u�V���|!���zK�}>�M�f��cC֜�c���b `^�T�]S��PJ
#�)�0&�	��MD`T���5ǉ���߿�nݚL�c�|՞8����z�3C��5<������4,HC��^,?:>��F%�����ibP8V\�>������φ"�X��/DGY��/y8m/�ࠔI�-z@8�C�KitwsMk���v=s�nO��)w��Q��{�Z����\*���4��K,��v7���b���hR���s�Ր�~���
��͌fH^�@�on�ʊ+�iG���}��t���@n/b��\q��r�lg�: r?>9�8Ux��Fo�s�:C�����g���1Zr'`|r<M���)�ÃR�jX6�,a��Ռ��}�
�١��OevC�㦧���֎�ؐ&�'����:0�#B���f��^�;�a��@�3봕u��Y��,���z�"����eۻ�i�%04^RnS[�t�t�U�JBz}{����ǏU_f���z�5��0������w=9�|�y���*�Sw�r���S�9�:#Q��I�]�e+��J�dcY������Ʒp��� Az6��S�Bp���4u���lej<=z��k��Ɣ[���C峿ψ=g�rQ���/��ON(p�9���̻2�0��#��l"g����i]g
JǛ������<7��ǐ���5���`7��t¹8ɐvn��1� ~.�`���w�qG��wY�9<2&ӗ��g3��^15��Y��UJ_��F)޳R+?���7����|����������W�qL��<Lg���J����{wo�	6N��o��]�N/���<9��"��S�5�a�g)JR^h��++^rٽߣ���q��dK��2#�1���jK;z$��v)��7XO��vѸKc��q��`�;E�٨�����NZ��v���GF�f��z����.s�²��,3Q/�V��I���n6x7��3f3O�J2��xK6--/Ky[��vKцonr-:�m{6�=,�8�$�s�9���+�ww��)�^J!�����+�2՟��q �g�f��g���p�f��=���0���;9g�#�ʦMW��S���:��t�-���������`p�@���1#�MzV۠���&G�rZH�	�hs��#?(Ӭ�>=9ߟ��ު2�O��Nz�Ȁ�y.��fL�;��?X�έp�<6�Ѷ��0���Z�S�}ux�>1�A',d 6i��9C��M=��!�����g��2�_��_S��O���^l�$��/�qH��!�r"�m��5��}��V�/J���Ab�Ҧ�斴�a�r�_���X�ܪa6���X{V"`c��b�5{�R�!&`x�MRL��)kn~ъª������xbz
���|��&r&,k^���a{�ͨ(�D#yҧ`2QD���FәB6�MM�yQ6�MQl�A�hnm�&���!�O�^��b�1�Si��d�� 爳��484,eS�(\��`��3n��(.�-�J�F陆�p�+
��	)�SJkR�������3l<A��]6�-Z�NM�w��}���+Vbzpb)W�.I��y�5�0��:����Mzy���Z=�s��-xm����O6Y�s�E���2D�a9�R��Ud�1���mN���fCwt��������-�~m�;����+��Mu�%'W<y2#�v>�[%���2w��M�&ǻ��?ğLS�����yJHD�ͳ>jQ~�}�#�uߒA)�#�`� Б�A��l���q�E�׿!xX����G�P�֚z����vٰxr��(�K����3�G(�O�>U~W����qҍ�a�/��H�S��)�Ј5��(�H����e� ���\�.X��@�Q�0���cĦqǻ�T�0P;�
?WM����=�r����u��ќT���U�#!&"��`��G�F��U�HZ��Ռݯ:ʭ�29.�A��͛ܯ�o͔���u����g��J0����}ʈ6��O�k���^�jjr*ݺu[�6����8C�ò���c��7^��'nY�r�ɬ�����8����O�[�U;S�KF�;��Λ���u;�!�K�&MJ�$�|�K֌J�>��|Z�m7N�giU��ٓg��aF6����E<��i�ౌlK�ɔ3�#�U�%���[�K� 3"�r�&)�M7P4Y���(ô�t P������62)aЈ�wՖ�|#�96�*:�}\N����A��Z����ξ�@�u�㓁X#˺Q�� (�M*�No�e���ƪ��5'�I��Y;ΜW�1�y�	2���nF��i�>y�¼RԢL�|S���·92lI���N.�|�ܢlR���3�Ki��j�&�ё��.�j)��ki�A���3{�����,�Q^�3��E�p� �����9���.�H�<��:�ZԾK���-�Á�=j+~�y��3����܃/(��[)|(������^'N+����`���E<b�����A~�<!�(�<����lc�p��x�!=o<E8�������a�:eM=�>Ӷ���)�i]��W��s���9%�c;2*T�9Q6����Kcw��ں���kK}�¸�P�<cS)�Y�	<�c�B0�:���Y����[BPQ(�sU�d������a)�*lF�$(U�ؽ�?0 ������3��nޚN�Rp9����[��>Ձ�N��O��\+�i&g*�klT�1�.��Vn|)\��cZ���q������Goǵ����z�f�(�F�[�nz�E�3o��޼���2��R�8�'t���%ۖ�&#X�A�n���v^�i��tf�U�z��a'��+f�ɝx`�V>f�/i�_TЌ���s�MF�ʹ���>1-�[N��ǰ�I؇R�ޥ^�z��]�ipxX�6��O��[.���	�M)}3i~n.��,��:#e�+��s��cN$|w���Ό�x��+%������a)�K(�� ���<	wo���H�Z��qW�%Ѡ|���;FY��޽5DbP�뻶�و���)nJH�J�=N\�����&�v)�z5���x�^�|���`oO�L�;B����l���N\M�/:�(������#w\)pU鄡��"�o��M5��]���6���:����|�����؟ƾo	�Oʔ3#	,�9���H���6��9�R��F|3-.��]�+.���=5�,i�8�v�.��p���z�[����q�)���%z�c���Ɠ ���q`�F�9��?����ul����u���f�p||B�vLujH����;�*�%�>�x�"]S;��z�L�/����5T 6��&#���@�&��eE�l7�����4՟��t�����x���$��e�vK�T�=կ������Sɂ=Ϝ1�@
#����A���ի����NoQR��`�I!�JFq��Ll6#s�GU)�d"
h4�Σ� ;� @�w�ӽTri{kϣ������T��f�NN%겲q/WϪ|�n�	�ܲ<��K��.Gn�c�����w��;�>�|����@���!��`��I��<:�N8���ݼHG��3����B6J�1�� ��2��߯�.�b]h7��Rr�-(�
6�0�q�L)�m�Rn%_�ԁf6�K��:�9��&�σ5�P���hp�g�����<cC�[Oҿ�m�I�za�x?�tVn/*���h=>>dś6�ֺ�d�s���n^�ld�g���)m�r˥+�H�z�g�2Ȁ��/p�G�&ލzH]�6đ��h@ߠ{QlÐP~���C���l}wv ~����+���<��v \��;̋��'��ܪ��Ɣ�.`6��M�"�"��2^�`!�����Љ�/"ﰫP��ʀjƯ�1�D�W���U��Rb$�l�PF�^A'"�)���c���Pn9ډ�%�J���9����>���[�z� I�JC�Uq9ʅSFN˔O�� ���ޚ�3 ӣ�;w Fp�0��)�]z�L�����SibbTi	����Fm(��溿�a+5� ��8*��CU���C5,j��^vq�t�lq�/��ITT�t ��L������2�(���Y�҃�(;�[��4ŐRnۚ��bP�}�`����������:)z[���6��<���(��#�G��9ڋ�/^�H/I�n�1�VVno�rۮ4�k�V�^ͼJ�k����ʨ�����+�9:E��.�&7����� Wg��#d�
�u����U�$}}.��i]�a�B��e�#��\H�jY��K琻�77h�}�"�KD�U��A��5�,M�r��s��E���g�ʒ�po:� �3�R.`>�K.D��0����<�d�:H��ϗy)��/��0��"]TB��&)��iF�!#�4q�H-��<k��M�HbC�o���5<+�I�Bo0|)~/�7��.���s��R��)x^�
�v.�F����Z�����,'H��&F���4n�}�K�8U���f��>}�$�n��Q�$	M��� �A�
�a����vN;d}��:����#��١���B� ��Mx12��N�V:�$��e���M�]wW��o{��ۺ8���hC���$�C�x�\���kz��q$#�ЍL[�Ncs+#���6Y�e9Gd�&?�F?Oߪ��rF��x���d��h�ٜ̦h�0���fN1��z���$	�MX/^H��]�A'�Qf�6޺=鋘�?�V�;%_8F�im�����Pe����1��1�2b���8���8���{@ȝ~F���Q7���9�Q�aJa��|�m�ݱl��A���f��m���چ�����x���hF/�Q�3�ʍebQ+O�}�G�'���<U�|P��v��,ɂ��7���X"���'�喥$Y��3e���Wʛ���A"�E�.qf��:(�� m%�_P����V2�3Z2�wP3(�l
n��s���L}�]�r(�L�"w�jin�'.�@�m��@�st�Qp��rK�Ȁ�`�;�7��~L�5�����[�V�ܪѶVNJNO�e"�hu|����z�A��=�.��
��e�.N�|?Z�{��8�BD��@l.��y9Ed���n4����zN֨�����U��E��OG���d�L�N)W]]m�Y�סƴ]�k�ؕ��!���qV�(�rbT�{�Qn�3H���[�&FND�f�^{҈�-�U����i��f�`�-�:0-ϐ<v���7ϔQ1��W�ܴ���������_��b*����z-�������6�v��4�^���VX��n]��W����{�^�v-��{�}�7��ι��{�BRU���H�"���w�B:|$��!T��涧���k�������?��<k��=�h$���9���=<<<<l�P�����++0­� �6�a���t�$�>��WK��{u�+*���E�$��j��t���V�X���4����0��$F��p<s;6��M3����[���L�)�N������3U�0"�r~�r��:9AC�AC�4��D�* �u4��D��r�-E��rܙcv����l��4��� �d�hA������b`������L?j�O�jHǇ�ism/��,y��س��{��F��<�_h@�$��
��%m�0�w�Q�n����s\�op�����ﳯ�罽��¹��ʜ���k�������������Y[p	�N�6/_��'���w���0P9v�sBq���>��]���:���&�a��qX=��n>pQ�v]��!2�^t��I\I��䙡C`b����{	n�_�x�������d]�P�5u���b1�4L?����D�3/Ex�K��&�W��}@S�s��כ��3U�����:��z�6G?�`�Jj	$ܢ>��!~+r<ܿͭ�߿�mXo��о���F���n�P����[p_/F-���nmq� ¨�lO��c�Q�����B_�x�PrGG�#Ա
� �X�2v�Q�b ��+�kg������#�b���1_��a����+����C�Ջ��X��Qy����haE�l���S��f[�׵�5'6������>��I<�\����=T��:�7��"K%R/�Z��E^�7�'��:n�vѸ��8�I�m3�m�k�F?�9�A�̜�6M9�'Y>�GE�YzV,ؠ�z��-ȧ�g�� FN�Ó苭o���!ܢr���K�(CC�W"��wt����"W�K�zf}Ul��fn���Nէ`�7������@"a�E_w�>jO��#�[8�@�)�A/A����<Óyu%�?���$��3���ܞ�� ᖕ�6˖�Ҳ'�gm�v��0tn��L3�F�3Sa��#i92�9�r:$e��D�i��,3��DEQ�ލj��{����4��+�䌘�k�w�٤�$T𤎾ٺ',ݢoD�"0����W*]Wf�lp�{�-��#��f|�`�emN[_۔���$�S�l����?�Is���%3c��i��"�=�� p�`,�-�g����j�����=�qD/zZG'��?O�{�$�w�!r�0�C+ས�dĉ(��;�WW�?���ʮ��ZXq9�D��"!�	�"X1�6	��fI��^z�Z���zZ]ۿgЀ�jn�Y���gy���ia~�'���/[��S4p�O0�Ɍ8�� ­,�0�Xa@�D`cF��`�W��a��k�!1c�e5,5*f�iГ�-3ߢ�r�Θ{ڇp�g��w��j#����	ud�eC:��8V�[3��4j�`ӛ|�8�clѷ�
�N�sB���(���w�0ws��M�I;�>���.~���mJ���T�E�c�`ρ�^�~I ;��Ox��M��5���@�G�3(� �s�oߝ:����gs�?q�\�9�}��~�aLB>���r�̻��`��R�������+�\���C�X��"%7����#:���^�08*��nf��Q�^7ǐon��c�ٶ����kQ�N^I��
ldZ�	���VWwz�
-�"���#~��9n�I��x�+���^�̛�C��|�`ڳy����r$��y�6q4++��g�wgv��%ء�P���5�*p*!	�	l?�O���ɥU���l��(�!v�'��{�����bƖ�̇�O������;ا��	���A�J�F��Ԩ�0{�]��͒�<1�����y	�Kn80؟&��ӳ����	-�-ěWW�ajWw''5(t�omk?m��ᶶN�[�e��������L&?����R��.Ӎ�s�VN�ES�F щ��,܊�#' D���PK�jS?СAJ��d�ZT�h��=���Z�ұp+|2s�5�]�­i�n�.��hc�菽J��=&T.�p��F�ǳ��I����ͺ��L�9ā�������[����j'�ACH�p�I�@�]�f���ؾ�����/._��u�����8�3����D�>tPy��_�Y�H�=�7�C�9�3j	�!��-3���έ��7 ���}JdO�
 Q@��h�1����F�d�,B�7@t��H�_��*�`r�y)>iS��1��NISY� �"����(�F�=���=1 6��m�	�<��><�K��˓o5�>R#�M�K�܃p1#P ����q/��>�0B��]UP���N��.ށ66S!�bV��}�4�?<���5�G�=S�rj5���7�/,l$��L˾B<��E������q�� z`���Bd&��2�JR~�%nr�}���X� ,vLSg�$����4/�|�#��8qL��W.�|jxyi��ۻ�y����p�#���P:�T2TS�NOH��p� "5���u����zs���y#�Oл;e=h�.��x0¦F��[�����U�V�ih�h/fZ�u���u-��o����#�'&���J�7é����3�����B�v���z�FCT�`��G貐1;�(���6�k3��Л�&��W�b��g��GbUO0c3j��D��rz|�=1�=8=�OO�p�[��T�ݓ69�T���zG|����dȩ�l*`_����`
��{\�|ҕx�}��ߑ�oq�ӯ\	.�)G�HNXU������.��9��+�yS�o�U������~�������`7����ӈ���rP�0����@Gʷ�����S�
E��|_����,r��	y�x�n�[.O�>�附>H���zmͥ&ܲ�\�K|j~�+=�}�BߛUe�	'����lV�'�ee�<�ޅ7�����!���|Ā�INy!ܒo�GV�BxayAX�afA��L�p�a9Fv_�C&x��:5�f���/��������f��+nm�Q��|Se|�v&m����������4�A����_y���vKk�``�뎏�G'�KݬziP�
VY%�V�����E�<̯b�,�O�A��)y�����έ�[T��	�� Db3����=�����C��3�[ÑiK �g�gd$p]fnq�?�ݘ�mo�Դ^��?��f���mܩ*�+=Sߨ�\X�m�p��ӣ<Z�)j	�x�6pB:�I��6�n_~
@^��&K[�Z�����/��}Ws�E��<����'�>��[��֫ؒ���͙[T��p.�p������j�z��"�*i1
�3��6�@�k<���70I���m� �W� /=	8һCE)	G��O ���>AS��D;6�u��AyY�L,�`�P� �0�%Aj��Gx��� ���2)ϻ�8�o]��D�Sl�aW#!1��� R���Ǖ{7*�"|Asd�y�,�Fpxņ�ä������n��$t[���+��2��Y[tO=C�%�`!��	�eo��.|��ru���:G��^��5j5�k7�01F��gcM=�-	�b�QK�L�D������V ��0����y�aY�i+� ���KO�~���� ��BfЫf�#ư�16,���ᰜ!��V+��`ر�#��B���T�r�i/�[Qf�U1�٣:�g��1	��,=F��t�����l��	`R~�o��p�[_|@o'�������t/�H������9����]6S+�O;f?G��$�,ت�hw�O�zz�J��%�_���������������$��+u>^6����(Lt�	�V�m#��  f������m�~��#/o>����8>�_�����g�w�[?n�E%T�O�f9�\�lTW���� ��=�!;4 ��-�Fծ�U/�j�֘�%�b/��o��`J3�!�y�a&����ے0�kD.p�~�W��~������}5]��\i��V}A�c���ʲ0B�k�c3����u�S��(��<#B:���BšSP��j�TxA�D�E�I"�KZ���"����I���ywR��$6@a*�U~��{�R�>T�hØ�.� ��f����Eu�Z�az?�*��V������h��p2�v��B��ښ���N��ϟ?���2N�G�ޛZ�=1��>�=��C-f��'���pu5d =��x.ף��k�|���X����v��H:������6���<KJ:�|O,�?�"'Z��)H	��Y��շ!d��$3/���7wQ��$��)���&�]_z�p�t���`�`h�� 0��e;��y��b����#�%܊�Xm98<T=Q'�'�OY.3ºh���)�.*�|z_ڦ.��0_q��x�q-8 wF�#�/㪴-L����º�	�!�.�J��d!�2 >+}�������ل���{�J1��2��8�(�;2�3�A�����РH<x��J�F� �SU��b�f;e&�X>��n��(dΙB�\9��Y�6��1p#��"��vF��M�4H�J�0��&�ã/�����e�$Gt�LhD� �LR8jx�ay�̰=tk�'�-*sI�
f�S������_��(����
9���.T'���ݹ��x������S�/fN0������>_Hy�נe}sj�]�*�J�hE|���l28������_�Lm�`'P���릋�Ьzeժ4DFf�=�ޙ* �cl_��95���K�={���?�K�ٓ����JB̸�|h�V��+�wc2�gE��~�3����;���b����ی�B:s�P����t$\,�a?�zD5�O�>Lϟ���id��u	c���7=����]\M�B�����ɖ��w�ͧ?��~�^��I�[�\�t0����W�}����&ĀH�&�3�n�8�]*�E�ұz>�v8��oJ��'�md�3Cm��iNSS�����Lx��m�`:�?H�iq~����k���E�|І��(�3S�e��O �M��cT�o�m8'���M��)�a�����Y�t�?�.��/�}I��#^��q3D�
g���7y�&���a[j���� kB�g{�;8� �������V:<b�(f�b��k�Lj�g�͑+ٻ\q��}R�<�
-���W`�Ue�Gz���6���{�)�OP��>K����S>����-=>���_�K�G?�/��N-j3�;'�����7�I�[��c	�UJT8KN��l��-����:d���6!�[�ňɩ��{]<�ۗ
#X���r)�u��䁾��%A�:�ʕ�"}����N	e��?6X�y���G�Q3`vpH�w���4�v%���:��|����7�<�����g���不�K�`��y?�z=�S�Z�[���ӓөI���-%��?:9�aHO�=:��w��׿y�����O��ª�2�[��a��.��֕z�{}R��B�yW�����*���R�g�����ј&Ǳ<3����H���S�p~
M1�<�A&��w៨�`�+���{B��}r�l@��M�|�����3�m��J�>=�K���3�Gg���_�W����Ե`a��/�g�ԏm�m�βi���42:�&��I쒰|��AG�#���8�D�k�v��x��5�hO��(Z
�(E�v�}�"Oio���n ����cԼ�;H�!� ��F��KT1�:8���>��;��p?�J���-���#�Z�����6����~�)��-�b'�G�;�p�$�^e���x�Tl �T�	r��/�X��3���dbTC|��I��Nwiᔣ�0�a�)K,�a�@B	�����?������O\��ĸ��O�t���Q����PQmG�c�>q;���kv������6;���b.fKLbǳ�[�{i[�1Ftj�����m��}vk���#�hO܃7�[��t��Φ�nx�c���5w<�˕���tؕ��;�]�IyK8�QA���	�RF��% ���/��y�yxP��c�T�A48hF�a�)#;L�����Ո���	[�s�C5��X!�����/�X��������5k Ѡ�4�o0CΦ�313h>�L)���p1��`*��2����cix�_��v1�v	�4B�铼�0���	�3z����]H�������c	�>$sD'��U��y�&�{�7�V�����7�_C�V>����KZ���LԸ�q冚����h���33=::���	?Qg|W�Ql<7tГG�`cK��3�}��8�|ɸ��<�>�x��'r�}�Cq>��Տ�f��΍1\��r�ui_�C��8O��(�*twvt%L�a�����ѣ�ill\�ث��?�l�Ĥ�}	`��p�P|(x��x9A���#��s|���N�v�,�q����.n����z���#fc1֒����}��T�Րp�/�~��p�-%���/���W�z#A�^1Vi�'���Mlr��$���'{@�{�_�fՓ6��P~����:�FY�ܝ��`��6QY�:՘x��x�k�=y���I��y��G0cC���W��Ⱥ[F�@O�.z�%̷�G�&4x��ʊ���.��c��A,'��p��+	�[in~E��e�x�ɕ|�7�(�����O9j.�rÁ"�I����a�������]���\��	�]�88�z����}���09�lh�Ʀ*�a`1�AѽMN,��pF��g�i����e2��mM�1�:99-_�]�������J���;t��ZP¾1�'�3�!g�0�Dհ�ġ��e�V}��h^����L�}u��ڢI��=2����Lq���[=�k�onĵ�O�8��v�Z�"��ч���+�C���Y�=��պ�$�S}��W�_������S	S{� ��2c��g?�3P��+���Ubֶ���a�����2i����0e� �TL�\B�92W2��/� ������н�t,��șk���Ų3�fF8;}џ�+Ȣ�oh��7�&|�j�{�_qh�L�33ɨ
��D�fQ0#ò��<cZ�%{Ml�v�329��,�3k�%r�D\g� |�ѐ�N���~����*�G9�G
�+��x+O�9�z�?/>����5�-�D��>ԃ�/���A
M�M��u��!�r�3vdٰhzQb��`�F�f��Kn��ba�$�����q�>���ǳ����^���xВ@a3zΨ��� ���+�TT���3��K�0}"ȲA����4L0>�[`5�C��Jq`�T3�����]v/礪ō����v��N	)Ouf,8�+��~�p��G<n"�F����)>��t���q믜&�G���U{�Max.�I1���'CP��KCb�]�s�
&�ؙ_̤!�	�Fg�+����!`�?p�����������^f�	����>����w?��G�ےnT��W0��d���	�!N'�>���@<&`�
'	b���\�v�;J?��ϴg� �M/\�2��u��|ke��f_��9F��;���?��k�♾�Š$a��B��{
%�a�M�̞1 Ʀ-jK�L6)�!rd��J���MC�#iBq��G%��Z��S���e�L���i�@Α����㢔�<�q�D_O�R[x��Qz��az��^��>�199� �ұ�~�����
l�O9�cP���	��Eo���w�P��`�CÅ�
Nڄ,��t�;v���/h��n�_$=؅���NAݒ�7���̒�,-������C�n#�Qd�mg�r�9pS|�U�����ǌ>3�4+쎮�������hz��U�ؼ�j�Y�hi>)K�B"��\ר��ډj
"��l�[�OF^9 h;����n��3	����g�*��3�m��5T�k�[��:��[oln��8���m_��G�b��<�][����a�w�)eӢ���e�W`GƇLH�Ϻ�Le��ǵ�m�~��"���U<�/����~K�tm 1���c�:ViX����fV T���n������(fAB�0��Yr���	)q�w%Jq�QNAo-�7Ɣ��Пr1��,�K(�Y���(ht�8rh���2��'��L9H?�ad�j��q����L�_�%	���`���g���@��9sa��}��o@�·������	��#\���,�pÞ��:�e��[��=�[h��%��p���2˫����;��|v��޿V\|�=i��N""Dà��d�'Rn���iP���^��3՗�8�Ȗ/���`�6���&�Q����7D�l*���O[�1˳���yb�G��Y�0vq�w��FǶ��ia[��f�&ȏqJ_�)eQ9��-� �)���%utaABzG_x��� �_�:��,�>'o`�E�ӳ�:EN��t�lB\]�Oss�iai�KdA?���g���\�|<�j\D!��7�� �Յ#'�3W}�kD�����qs�S�P��VgҢ�{�d��
F��N�/��ؖ�L�e��G�y�tZ|Ŏ���]��\��w�����f~w��ʷjƋ�*W�?���>���^ԇ�ρ�>������Tz�&�5�l �,���m�m	F�f�n��H�FL&��+~\������R�(�a��<�)^��p�w�ᖾ�]���הS��b����A�n�m�f��3ec(+1�N�c��Z�G��6���d&��A��D|�h�j�lD
>ϑ��4Cex6�
u��c����;9.a��}	�j�$����>`b�x���5���3����t��#�C���vZB����̻�J��/���螛Z��.A���a�(o�:Cjܟ��u'm힤��L�%���DT&l0Q	��K}����RO���f���A�����ꏟ�"$�!�Y[�n9zwx������qh�WU�-���+}���Va�{���G�V�r�a	��Y�+�;��\�7<u/y��sf��=s땃���#AU��T�ԷiP N���`���w�3�}�n%�2(�fB��i��� 	�� �f����U^�^j�?�]����Wښ[U~�ύ�n��;�B���w!ᖮ��Nh��[t���P��2��[����-�TY,�����[�e��d,@ ��  �����5`���^�2�Ҳ@g�_�eN2�R�'B�-}�e-YJ����K��'V��W�`@�9���h��V,G���2t�ǌ3���=���VDc乜*�� N0���+�oH����i�_01�qs�����;LC�����1q"Wثe9�4��g6���T�� P�8n�2��x��S��)P��׻�� pJ����rE���3���D�`)ء�"0��J��K���LB�FgW�I�q#B��Njc���l�������p2O����&����4�~�����̧w��Wt]N��-&��,,l��s��J�O�/��ԥ��ʹ���	S�;iU
3aM�/�k��������>TyfY.B�Ħ�����������y�9������z�G�qQ���V�w$��	ƀ��*	0Y5|���:p xՋm�q�~�׽��ֿ=eQ�2�+��?��ZB��9�Gt;�7�X����9�[��#V-�57�i~n�~yy�8�zg06@!o��y�G>�ȿ�"�p�o��n����Z��r������7�����r��
���C�]�V�������Ի;T��8�=��d��|��WV7���O��?8���zc%�����B<���<�ӧ��˸z������i�F����TU�3=����?�G��sX�1�+q�����H�ȅp�*��U��/t�Ǹ/4�����B�@�8�����+��،��d���>��?��^�%��I����Nc��r����l�K R[i��ٹ6�9�7P����4�=5ɗ:!?���봦A23����y�m�&}.~|�p�_���,�)��O=9���[�k�b��#�9j��<t�݂���j�k�͔�~�W�Zm ��c�@�-�aؓ�� �,���J�1Pf��*��^0�y��g<7[�cbb$=|p���k�>N�e�-����{Vb�0�]�2�F�G��21�kޫ?������Jس��Dɩ�������4���Mn�ˤ\��V��E����'�1s۪���[��̠D[X^:ЕC��O�*\���;)�=��J��O�+�3���>׍��/ך������U���7T�d����a�+�8������+�e�G�3����v��/I��0�9��bdPD%�Rxe�;'N�d&a`ff!J�)�*ʰ�$T����_ FGRVdF�E��a;T���&R(>\n�a+^��FڵQT���wޠE#�����z�R(�u��>r�<"2�J�#8*7�Q&�	���#x(},�I�����B�� n�lȱ��.��=i�"��Z%��-iF�[�ˡ�����ϛb�ёj�/�0��k���^yziE�H1�p\E�r� \l\:n)��(�5���E�id���r��-�	j7�,��c	C~U�ڶ�®;@���M��wXb�K�{����|�P��h]x\0
�/�}�
ox����@ЯF�zǶzW$�b
m}-���B����m�����챭z`�ۚr�Yb���4TZ0�-���W~�L���.N8u[���L��:�`N�L����De��Z_���Md&��r�y������������Kv�{ؘf'��Y��شJ�->t�Sη����7��^w��O������x��G�o��^p%����S}����X��[lჟs��V�{9���3��]��uu�hh��uF�|�tU�`^h�{xm�D;�����q�ga��t�Xŭ�+��u��|k勰������G$u���E��]DC=�26�a����g���L>�#.WT����Ķ|�m�/�&`7ذ���Yo�Q��q�3s�
Fo�-`���@�-S~@ e��g��~���l|���Ⱦ�(å���jWl0��@?,�h��l�"�,*X�@ev�0%J\N~�0�5��=r��8����޿_�-��/N�t
Y�A�Z��\A5W�X��&h~2�x��F[�P��p&	����(,6��>�	e�����Q��;U�$�ȓr�.�@�	���<�� Юr���ux�o1��	)��.哣O�g*�ږ����g�������=8؝�&��Q#�J#GVia�Ki@_��n �J�eƹS�-�&�������_��o��θ�/8��k��9�K���1�S������S�\�o��0�
p
�Q">�k���m�l��ŉ�0,Ċ��tR�,��������zI�W�ްv[)�)Y��-�Lw:O�A���B��̤g������U�9;r�R�!D���7�\����G3w8�1S������ ~�t�Q�C)h~�/v�#�+�(� V�<?��F����0_��Fiᶒ�#1�C�G�r����4jJׄ�UV	%�s#�+�I��g
3 U'n`��ɸ���_5
:��Jй�Cb�'"�#b�\��3��\+������K��\O���*�
����˘�:�pK���?��W�
t�k�6<��N��P'6����.u�t��*�bF���_�%Q�*Mӂ<����F2v�B� p�^)K�:����|�D�{�8x�F�L
��:=V��dĐ��GC���Ki�s�ѻ�(�;y�N4n6ܑ����YL�Ӊ<�q�EtF�1������`�F���c`3K%$���U70m���8\I�_� 8���JlJ<�����%&��UF: ���[$�^]����c]� i�j$0�HR��/�Lifȳ���e�/�\\�f�6w3�mG����=���8�����Xʖ���Tūs%�zw�)�"mfC�����̗��JFݧ���M:U�ژ�;9oO���*/ڕ��`U�AVГk����tճ�m�����9���"A�H1i��r]�r(*��4�߻
7���/^Ŧ߹8J}}�����t��H�7=�F$0twr�_��
ࢯ�h�ܑ �� �>�A��m1������Rz�vуg���Nkcs�fh*�:m#�vJ��Kw'�ҳ���Ȁ�!	<-�_�>���'�a�/|���0���E̲ί�ￛIs�VW�8E��C�eC����x�~O�pX��h�ɠԛ$�ʈ���>�]a��=
�p^\�<Qn~�+���KP�����sQo��"�NJ::�R'z���-�X�89:L;�iog3������t�����埤{w'�-�cJg�prk����U��|��4ln�$N����iaq5qPB���a[\U/�R騍���j'n�y�_�D����X�ɞxݕ-��ٓ���Ez��t��P�ϵ4IPW� ?:8J�K+���r�U=����ٳ�?0�~{w��G�*G�-M�{��e��J�	�qX���K�[�ݶ��W�8f��|#��,|�m8�S6��6�䑶���?8���NKؗ��gx���N:><�<�����A	��$<2�R]}�?�C�3o����UP:�hQ(���D�j�o� ��G����f�� !,!��)q-�����l�uA��GMfp0�`�F�;�|]�����
�1�|�8\����9\��$`A ���t�r�Օ-�����#�����z.L��@��6�u<�\��(^0n�7�%ʉ���R0�h7��;{0 �A(4�'^�U�����.�;R4XjꋤJ�6	�B'CK����$���;���ǿ�u!��[�W�<�w��wy�9�Jz�L��s��@n��R�Mw0����V��\�M�֔�q��'s����_6.��I�3�Aq�?:e�F��FC�[!3+��cvxNdSI64��טœp��0bfD�/屘U�2KeS�9�h?AC*�q����v--�*S�DF��mb�J߸��zaR���c��Ҕ+�~ �{_n%�h�-����t�O����\I��G�E����W�S�\]���^'*ӕ́��Q��tq|x��ONWQh�פ�؀Ӱ:3�S�K=���;���R�rQ"���'��)�?p������a��=�4�F¤Q������Wn9��v'�4"�Fթ;���NmG�G;Ɗ�m[k��kN'X���-K��}M+�.�]o�Ae���<�/qO8�����B�q���+����͛�o�
�W(�N����< �Ez�H(��NM{ʂ���١����F9:��f��z������Je�<�c���o�Ҥm3cʠ�zV��V���
�Ā�v�� ��a�6C߆�D�z:;Ґ�ˉ����ە�d86ue �l9�Ī^�oo֥��xlw���G�"t���#��ūNN%#��0��|���_NL;��K<T�ʒ<y"l0�=�;�[IP���F�\��U�q�o V��%���{{�:6�nQ�H��[��0��H߽KK�i}u9���M�'�0��0��JPRy���{�~l+,�����C;��im}#��/Y��B�S����n�w[ݑAv�76�T��X����U��:�[	�'{n/��@��Z	��Ez���ﳥհ�[�%�7/BE��˗i� �[6>y�̛���n���⒄�m����sܟ�j����I�hl��E`=��Y�S�իP]�(��Uu�o��,÷�1-1�l��`O����7Ar�tu!���lk���R�0�}�L�V�;����r������,���e �@��#�f0:b ��!Õ�F��O�.�2e�#�
!fŔr^� �g�!��:�<�y�T�	F*Aգ��*}����JX�5Xy#���%�E�
�L�C��0��o��|().~�A��Oys�pD�0h�QI��Ms2��L]&��I��G��<�X*�(��3a� �4=p@̤��+�_��b8e=�ޔ�6�y�y��OAT�ⓨ�M\���k=\O\�?i3`��!d�F�!��)��s��"��-p�3����}бW��H�4��M���]\I��W�0<�wV�����@!������h�_��̽&�zFq����F.~�Y��ݪ� Ov�`N�k�W��;�&k	���� �ۈ��Qybc�����+��<��
'�.�� ~���a\���V0� @�s~r�6r�:���Hwz�p"t��&�m�������`�0a��ͮ�(���#�|	�!��.�W7+`�{��{|��W"�6x���O�)�P �O͕�U��(��y+�RL���?�Qq�5�4�e)��/<:pt&�꼛������w��wذy�g:�.	W�V�:����L"Y��I�n�ڂ:1�,r��}��6lp����\�!�"�~V
DU��4�=<���`�Y�K	aཪ�Ieg�2�7r2.���Du3�ۀ9x���Ux�Ȿ�N&��X�8�'e��T|�_~2|��h��&�[�G��Ŭ$�&�-�B�U�t�c%4T��R��p������0"l�I;��#m�vuƠ\�s�1&���@�/b���#]���%L�RV�
os񀅫.�yN�W"	Z��W�я�9���DBb��:K}}������XB��5@H��~my%��g�H�}�]�y���2s;9>���<3��l�n�h���QOF�LG,���(ەh�Z����.�=��ٌ8�k�2f�.���8�xGx̊��x���P�ok�p�&�v2��}��?ǂC�4&l��+��	���!ܲ����)fn��~�Q��=	��;[O�[A�G�l�T����e�Mg�X����ܶ����$V�%>}0,_?���h�<G���N�8*	�#��޽{���&T�v����ѱȅ?[SwO��i�鐉-��������s�N"��i��$!>	bF�S�z��9'�.�@AD%�1�8=[`R�������;wL"~�-~��������W�p�c����8�ď�� ��<�oή��w8'X�)���U-]�^y��j��\R����z$n��'��">wt l*@He&-f� 3��>�-EY�-�JƩ!�w|Y:��Kx�#��8�}�R�EE���D����l\�G��+��xt-��.e�&\)C�5���E�������N��}�*�pf�!��㨵8м�0'i�|��nw0+d�k�G�	�x�-���w㋶K��������b�])��	|� ����R���8�<�өQ.ݛ�A�Nf
��J'g|�_�x�����������Oӳ�����M��h4߇}ζv��h��,�Yj�gP�f8�%�«��Z%>�n����էw���ou%�O���*�O�a���\y�?W�v��m��`7���:�v	K����p�6����t����ie]��SbC2����f]�=!�O"���'�B��	��Lh��%l��y�U�P�� >������\v��K	�V��,L�G���:�:M�SՇ.3aL X�S�n���#[P���	���Q:@ٞ���DL6X�s�-�#�G�q%G����^�C �����N�!�j��*;+M���-vr�1|�|�s=��+�����ǲʑi��K1z�%��}7�J��X�A��=�O���]YQ��
�#L|�D���e��CfLQ8Ӂ�s���q�p�#���B�X&140��:>>hkϞ>�满�E�L��ik�s�����Q[�`C��Al�H(�U�c_]��ѡp�-��Ii|�4�T�ď���So_�gL�!�Q�������/����`��M��%�	�x�$oupB�`��ظm|c��]�p�۠�����B���%6�:�86�q,3����j���\:��u�?�E}P7�O���/ם/r�W��z�7��Cw�A,SDy�=���^H���a�*�2/3�,�p��/�8���'���mK�E���'l���H�L����@����5:[�F�R �p�D�Wf��{��A��]!�|����� �������y��<�$yVӋp]QD�^D��H0��:Kr��� �o8>��
"2Ό+�¬��0��+τS�`�8Ne�����t�9�7��3@�9F��B���6��J�rƣ�l��f��
��s#�0��|�K��g��w������ڵ�Ʒ���{ӗ_����+,�[�L,��3QC GqE�����p�S�"��f�?�@��Xm�ơ1�m��"8���`k�����P�h*�Z��H���Qf�����8��S����O�C��B��~�%��~%��i�B��4a����j�k���3;F}�S���7ХQ�X���G�&Ұ:���^y��P�h����a��=I��s~�������]�p��g�U�ӊ8�R�b����n�[]G}
�{���oKX���J-������+�&v`��~l�>~�(}�嗺>Icc�D;��i�(�Ix+vn�Q�� �I��i*C�S��2u�F���͏�m�*S�#�p�hS�m��G����ɣ�q	-�SqLs�R��g�[� q��c��{](��DKy�|J(���(��l8Ś��镄A�Fh>�5���qBir��7坯x�5
�~�Ȟ��l0�Q�z�M����}O	�~���C�P7���Y�w��dV�B���P3
�͇�Ee7<��*K��11��]�9f�Cy����ʟ��B�@DE�1���$\|}:���V	��ij�X��f��������678Q�H|�˃��A�f�ٰ�0�,!��� `T�ZS�X�6^��K������^��(L���v����N��ò˞ҥo�ޡ[�%}��Ŀ�����jU���'���p��C��.���������cX��G�����	ꎍ�x[����$ġ�Wx���ؖ�����"��W���B�����6N@-��3���t�ַ��-�٬T �{���Ω�B{���7B��)�G���Z��`��)�������U�A~��74��iB42���w�͹
>���NY�Dl�����*}����zY��Q��*̅�2G�H���.�Ǩ/���3��D$Z
��G":���Fm��2��;���RphD�;���7���pL�����e9lc��,��!��	�q���xAd����l�/������)eF<f��:"���LM}�g��<��@ �u_]	&�����o'�p��_0a�!c�a�Y�*,��lTF�~rY��mw#L���2�G�c�{^�N	�������M�t��?T�ُ��˓�5C��
�u�Y�.��q_{�W����^��ᏻO9�����f��J\�s�_d��}]��t��af�Y��ag�#9�ۢU��)�O��?��4�?�����3\-��A{��������42��w�/�@�э��P'�Y����dO[��*z���W��@��zѿ)؀��K[+|&{��ׇ��Bo��+`h��P�CO4%VR0��U��4{	u��3K��U&N�b�+h!����^�g���]�/;��<1��QE�A`��E�����-$H�y	s���"І�s��uiO��x�|_�}�޹�h���ਫ਼��-+KQ�\��"�H�N��+q�/�!�D �7�c��;�	!qL�`5/�"5Z�����^p��]p14<b!�&�$��3��'�q��А혚�J�����aN�$m������Ц4peK=�Ve��S�I�&�?�O�>J���!e�m`̓v�`�l.��[z� ��{`"�ʁ'�1�Us�h��9:g��{�������r!��l�ǹ����Mp�o*�3����+���왱��S+y�e��+D���Չf�x�w�1 V'�t�f"zOVn���p��ȋ@k.�1�<�YxI�A-�3��Gj�����|�P�=;A	�W���]_�K�0�`� B2B��6�*%H���J�i��/ވ�=q�0)|�klw�i@`�pz�.�#��v��9TC^�3��{�li�)�L��F��F�����JE�"f�ՈB�����|�Jy����[X�	�uIق]v���e���;5$���ڔ����w:�:��/�b�#z{}�w9ie_����/uE �a���%Z����r�Ӯ}����:����{:M�0�A;��0���K)�n]^���;:��J�t"n3t8��|2�Ł:҉�#����[� D��K<:a���*=z���AV��x��1Kq˗��Ƌ*M��^���tx��r̨y�[N��`������I�E="ఌ�I���a>6w! 1�L!3\��t���Tkn#\�"J�%o`%L����g��C��.�Af�#����^#B,t��)@�B�u�"�2�+�N����c����h��Ȗ�h������AϾ���6�oj�2@���g��3_VXuu���x��".(F�K&���Gs#��F{a��M�#�p�QFpcc`�Xgp�r��Q�F}�F3\�D�*�L�x�Z|~gN���x_J~۹n���+���h�ԟ�_�"��M5����Qϊ����+����N�͚��JO�<I_~���ӟ��W&�>{f�wt|��.Gc���{��}��O�>M=JS�Sl��F�!f�Q�����&=�2l�S�pBn���n(O<�y�W�|��`)C��+���_>)M������ ��r��s������4ԡ|5��͖{�
,e	��a��l=8>T:�1�i@0t�
�惨�\]�\XZ>�� N��WP�M 3�L�f|�k%�'��_kQ��S�J�媊�;�ˍ�ԁ&̇��z"���R�4�j!����O��÷�^��{�kk���gw�ome����2�l0�������f�(�<�\VE�p|�)����M��ӊ�k偿R���rmj�Ryi,��<UJKB|����7J`Fpn>���A1�&��Gx�,l�/_~��k!�R���|�K}W|D'�����,_fA'�h�����<�� �Ȅ�3�w�Z��<կkЗ��.5��r|<��% G?����zG@��%����v��������+ߔ?\|��^�
8�ϥ�Gx����#.ǣ��N>_~��`�����'�mn{:L�D�g��^B�B�t���Z)�Ic�{~~9�~�>�|9����U����fgg����8"������H��w?�eܻ}�>�^NN����NZ��ϾOo߾I333����	I�%��DU�~5���|��ӄN��?ŵ7�;����W\!�h�Zh��3::xM5��[�x�_}P�c�A
āO�^B��r���Дk�x���>���O��/]˄�A�̔=�J��sr�.�#<|��?�7��lx�R�St��g�G�<�������&pz �t��_�=�kL*�G.W��30����x,�N�*����*�~�����e��R��l\���p8�|Ba���64ܟ&&F%�N���^���)	���i`���4����X��J���i||2KV�P������e�[�٤�2 #������ª'�,����l\�L��}(����zDHg0�!8Բ,�f~�|
�U��	?G~�w8�\]�v������m!�l涞wT��%�����_r��v:�� �44c���s����w��QAP��Bؗ��IP0<c[G���e��}~�Ƿ�YE��`{��NSWw{�bw�F0�TВ�;0���x���Y��c��шX��2v(Z�?eY@06�cB�7��p�Kn��-��ĥ���l���<(�y��^y�[�}���lFb��7�L,90�f&T\avEx����x�������qaz.��A5��{d,o3L��=qc�u��]�2�k�޲�O&_E,`.p���;R	h�K���t��x*�6:�����0����(�F~�'�t���'<�!͚���U*0`ݙ��t�gS5��}����2Lf�K��W�dn_����=�9zv����`�n��������ˮ
SdG(�ǋB�]Π��3�&����c0Fy��c��*3H��奅�������ߧׯ$ܾ{�VWVҞOBuG߸�(k.�/�>�������7Agq�]�[�n\~��dڷݭto_�� �z�p���Vpyt��?p>v���(��)���/jp1'?��VG[���X��lhR�ۆ��F�ޭ���@>��	���w��U��[0ȴC|`�L���x���E���y����*������M�#e���gŴ�a$u�^��2;���>��	;Hi�Uv�e�����У^�'x�C_�0t���78�|��X	���^-���U�^5A8��k�\�]�%M������E������l�)�n��kH��)������Crz��zW��gՋ����,\�\��k	�6�5>6�&'F��O�nm�o�� �9����_<N�C�߫��i��ة�e�~s*j	��l��͔��bC���jz���њ�=�*��f��һwK�̊ B*��T:V��ӫf`Ydp�G������㟙ńN�*��@!�HK𸸌��P�@���z��&+��>|U�z�P��@3�Fh�[.h�C��Y�ru��C���I}��+�{��=���Q������7��s�yo(�B�l&�����.�l�l�����Ց"r|塮$���*@3tnk�q� 1����ŧ�H�ff�È�����E��e���8"@�[�K�E�lkkb���ȀwWON�����+��Hv9r�s~��D胜�=�g%������+ߗ:�;[��1�R1�c&@��1�fѢ���rǊ�(���^�����5�3�
�����u������^vS�+���骆��L @8�|�����FD�:�;�)�	�fX����RW��Q`H&,?���Err��V>��\���vJ*�ƍ�]y}���$a�0�`�P�-�L�8����A�7}�+|�+pEH����=Wʊ+t"��R'N��'穀⽢�"�£,�#D�mt����TQ�������Ү����5��M\�N��5T�a�Wy=ؗ��>EetBt��W�p(��y����Z�]��������Nj3���x3Kqev��+��� �t����Êˏ���G��)A��}���\�V�M�J�+W�5|q�U���Y�N�Zzx��AV<3�Ȭ�{r|�r�6377����n��c7�i:��V�;lb�w���� �QѨR���P�����(L��v��g��� ����)�\.����-�AG���&�F�����G���5O�o��M��Ç�Dv�a�'a�+��� ܑ��*_|��_�/�g����s8��.��>�L�	>͑o5c���!�f��>�&����� ���ҍ�������(��{?�\�q������rW]o�;������\_H��rxè��A����cJcg{7��p����NNά����}oe<��m��rldf�%�utH��T�[�4�bź��s���7j;6Յ��ёa�#�Ȗ�6���%[K� �X�A��sRYN�緵7I��Lc���9��M�Cܨkp�\��`���,Nh��4�o�BVʰ@s�}p	����=P�v����'���;�Q��o__O��Z�V�r��z��g�i#��!���F;e � �v�)��0�kI�o�;��?��
^�H�#Q&'S�0��QA����KfkYB�� \�(��e
En�d�ٰ��,�э��Sめ����^ٻ1�ab���d�a��������xz��Qz��ό��7�M���;=5����\�hO�w����FL��69�������V�u�d�ȣ�`�fVE�Í�!\H�>;;�����)���ң�w���S����&Ҕ<�����w+�~w2��3a���1!�3��=9:f]��(�(��՟�P�::�Z��W�En�Y�4]ԣ�����E��$-oL��K0��	�xg�-qn`O^���8 ˝�"*�O�Y��N��Q�?� �N!�T��i˼D ��K�yo�^��c���T��2s�s����t����.a���R�F{�,���P�����bv���˝����(�e�,~��N�Ww�.�����T��'fTj��	|�W���ݮ��/a\5��(�W�}��W^����H��
M�c�GW�Q��B�v\&y�#r˰q�ǽ����4�Gb�Qz_�r�W}�C\�;.q�pQ����V�����o�I���yuF��^�E��As6ԯ��%W�yE�h�m������̆&Q��n�]%宺���F����Su���r�3�i��ޑ�b�芍�(�2���X�
�%��f��)�K��_�ƴC�9l�f����ٻ�Φ$��"ܴ"P���UC�/�͒VBŇL�JGWA�4�a2��4ɍ"�toOy�)�c���������r|�t�{�l^˳˄�%>ၯ�W�qS���]G�}ݕ�|��ǥ����q���H<�=�H<7���OT��e�5�,܎��@Ow���N���K����ڪd��C��N�OK@ꖐ��w��9f�b�^E�<5�W�ܒ�,�1���in~1�̼��U�8M��I�n;�iey3�ϯ���C�@��'��Z�z�C(�4�frnh���N	����qԯ눺T�1���-�3��aC&���(�0P<>����\A�P��(�Bq�Kĵ����k�rN/̏���CC�W�+��S�u�lO��ϧ�aL/,��K���r�1���&�����x����W_!宮���C��`bn��83>�t{6I!L����@ D��t�n�4��ݰ�W�^�g!h��x0qS��DGT0���G���$�>��`�0ݗ ����P�gB�9��/���!=3��9��#CihdPh��d����<l�/βg��ir�=X ([E���p.��F�����}	��c�mȳ��?�w���+<���>&f�Gt���ݨ�F�qvw�(�ƴ�vO��$ W���/�0�+��9=����>�<�A֕TG�z�>��0^Сa�z&5�A]:��! �a�y�t'_��6yvz|+[�� ':?6(!��'̶UW�=�
�/-�[�.H/�e�%7��~�'�"�n�̃���H���/��e<�J�cع��>����U�5��ݘ3^숣Ky�Ώ�Ѹ����ca�n�22��m�qD)��\�#W�l�nu5����9����/�dhp��0q60���AP!�,q%�|	g��*-RW�	��(�I������.x��p9J�Y��_��(�ԧ;���r�{�V�r43�M���3�c����S�L|s�eӑ404��z�S���+�!q����&rds�U�:�jC�z��Q{S��Oc@}�*׺�Ai��e�*��n#i���Y��S�8�{�%��``:�G\�K��U⏢�>x�������x�K�8?=V��e}�7��'��b@�x�IΑ\*�W`$���wc��ThXĻx&q���c�����ӏa�>��E�f����|%�]~gH�E�w`=_�Qkq���ċ��#��+��s	N�����Z�P�I�n�
�P�wn��Y��V��`X�7������{`��ܣj���9	��g�\C�TB*�������|��[�a	�itD����<3�ic}W�nW�$3\*C�Y�l�\���J����ݚ�%�v���v�f����J�}l����u�Oڗ�;�����w~�W�8!�����у,���������W���
�@��CC5:������CΣcF��~�
ȵ�A������3C����1�*g��2��щ�p75���쿑p{���7m|�H)�̗G�\���"�P������N$��늴���[Q]�cncVF��{�&调9y���4"�[��A-F�!` p�����	��tz�����S=a�C#���#��W#�=��@4�;:�R����M�v���^�z�0'�y���ű��fX0+���P�Q����QjiN&Ա�A	ܓijrT�O�@����Z�Fi}��x�*K#�a}zf4�3�1�r|�VW��`���>�W��@T���/��zCb6�hHD��B��[�Uħ+�104�����́E�-)��"�9Q����W��k���@���{�N����V�Q�%;�1�F]��s��N�+pP����#�a3~����2xbF
sG���,��5q�Q	��+�2�c:�'�g�n�ʂ	��-tDXx`�ʆ:1�&!h0�U��?%l���
�q�Q�r=�/r��\�7��},W��r�	&/Ҋ<�9>(uT�E�*��r^_�j�V-zp�n������Ϟ�gO�h`8����R[k�:��=���f��P�2_�x��ጏ����AZJ��wG�Zzw���(%��>H�v^u���	�C�^��b#R��������gϟ��<=|�4��(�I@�LM����榮�w4�c��%W��d�(�/x��ںxU��� �����_y�g��k� �TPU7zg�=z0H�ڱq��^�7�1�/| +"�!�N�(��yU���纞����]�C�S}<%w���WqQ%c2�܃:/q[y�7��qʡ��?B4Bw��Q�	~O)�l������+���s��e�Gg��[����:^�7��v�øć��~��{���8W�~��C���u�w:E��O����0&��:�n�]�#����O��֏e�aG���V�W%���E�/����f��ٕ���I�r������崠4��]�_J������5���	y&�Mckk�iyi#�/���L��7�ۢ�� �������"��rvo��FB�K�T�#���͋><�l��d��X�`�<���u�$4o�!���T��z)��˯L7s7>%έx�=tA�`1�\nQ�@�g�Ŭ����-�l&8%ܒ���y:<8Ԡd75���^�,hE���t6��5��MT4�wcF�3�=V���I�(s<��%n�f+����e$Maj�'C(�����J�AW����TN�@��c��$ԲLѪwl�h�m��1�zn�nW�[%|�HX��4�zG�X&M1�g�%l�3�w&x�=f��'�MmW��{}��x/a��tI�|"_y��`�h�̻ �Fy\9-��C°k/�}��HE�+M��$Z3!|qo�	��E��%�b.rTm��ޙn� u)��h���U�̀<+BÒ0��xϖ�k���l� ���f�K��M���:�w4�4i�׬A�袧E��zV���uk����b��l���b�I7��v��d`��EK�t���F��先�t��,hQ^��̱��֦�ֵ�E����Nx,j�E'����穩�Bߠ����%t�a
a��K{1�
���\-���ڿ�á6������[Qe�Cgd�q���顄�gϞ���?����q��Ps���R]?ဥ�`g��������N�ǀ-<P���r���t�L�����嗟���iz��#�F�����#�6�W@
���R����<4�QG��C 6(��Rgyxī�+8��X���G����*����<�4��"��]���k6-�qm"ܖj�j��-X�Q\���Fx�x~s��Ӹ�CXhp_������>�֑U��s(�ZV��Е�xuep_� �Ti��Y�+&-�N�.��Sy�%���2��l�%���n�������Z���������%CO����S.��1��xW��$�;_�%�S��Tl�6����\z���-�|�����7ߥo�{�^�z�f޽� kՃٹ�����|��w�;]_�;�m��7���ʲ�i�dp�mv�_n��0~T��B��&L�i=Š%B)��[�cZ`rC���8������5�^��K�F�C�c��xis aٯ ��<���Jr�9d�C���Px�|��=���� R�>�<j�	d6ձw�����o�B!zu��B�H��b�}�
�
vS���?Ė�͢S�s��F�؉e&���BU�JUx%�X�!T!���7I���̌Oㆢ?�����
�t��'G�=�/ML��!�|:% ����e��=M��I��9*R�3��H�_v9������ks�~c}'-�-�%��VVV��ޞ�a���QN1I	���]n1�%&��Z�6���<"QO�N�_�9�I�-���T;0��´�#������T�=�kqqS�l�G>�{:��ą�I`�A��4|һ1s��/lXݱ�a����Q*�Wu$0L׵�X�Q�ʊg����^�<���U�%�ʹ��;0B��
ϱ�(��x.:�#�a�������J���ty�1��w�<�5��:TG̊��ԙ:uߙs{\eg�!�Z�W�����	�(�,e0+^��^�x5���@ߎՋ���*��R<�j꟱��P�=X�b�
��L���l>�W�
i}r��0-�U��x�(����pu��m�A�s)�%���ޑ������|F���r�:jAc֝�
OW':VI4�&	Tq�t��-�E��4�ɻ䑟u�O�+�w�G�:�3=����p�Y�䁯K�x>��r9J���p�ҿ�W����X�(�8�Y���6�`mftt8ݽ;�?yj��m���U��u����C�=�*%��S�n/��]>ؿ0(��?|�ӕ���X��<���`�$�G!=�B��|\��W���}�P�l&X�9� ���̢���oww��o`�|��E��Q�a��o�Cm3��3Pn51?=��FA��!�O���bx�J@���>�A~�_�<+~"���L&����0��Wvt�������s��3l�j�5<߼\�P_Ɨ<����w ���k�\�0L��<����z�r��8>��~�Kx>��0~p�����3��rʱ�����.x斾�@�uq(Apsk+�m�ە�t`����?�O��[i[~k[�w����+޳�+�唏��w��y_*� ��>yyy+-̯�[,H>�m��*��g6�������3q�>��MϢ#|� k�ʮ�����cy߶��I�7�S��b��.VTU�$�d��s*��X]�v��\�~���S"�7��>�7��`ˌ-��:{z�Vl!A|�jj�>TC}23��ꗡ/۝,�l����t��޼^\�L?������]Z[ݒp�mXfA�HX<1{J�(0 !��*��jÙ	3.�?�4b3���f� $��-4Q*�U�$&�zG�CЄ�А���r�P�(1v������\��F�W�iZB���_J?����Ѩ��3]�_K�=L+��D\�L0s3r" �z��+�@��B�1��+�jg�P�b9��	�y�?��800���c}��2�B�a	A���=MM����XV�L�����6zlh A����)ӉC�`��s:Bf���Е�ά�?��o�/�:�y�^����H�Ӧ���+��T� v9[y^D_NP7*;i2(�x9�R�[��rX����3�>��ʈK'�r���ȢY)	jN�i�ghE�{�
�}p��P��� +a�b4]¡���Jd�p���)�R�֫ ���<ˬ�/���c�N�CN�d*K�ڋ��2kM��-���0[ڔ:Iw���{�1B{���M��t��vЦ�a�&v����މ����JLШ-y��p�[R�N�ΰ*rt���_}�x���A;U��Ʒ�	��4�r�k�SKK�|�?+)|~��B�hi�� խ��dz�p:=}r/���C���K�KK�����%ݳk��P� p��t�<s>g��Av�3�=ڂ-���+��Ox.%�B�Q�Z���������
X�9��V���n�cCN��Q�S���?��h�VZ��a�H*,�LOO�����?��g�Y>l�]-,������g�w/�Z���y�B�t���Ѩ��኶�2M"���̭f��(��]��o)�J�E�ˎW�z#~��B�k�����H�����7��D/�F�����z��*O���[�փWȃKy�xLE�4��Tl�Yy[�W�¨��ޱ	igG���Q:P��h^���\HW�Spڛ���g29@�DJ��nS���>:��\ś�v���K����C��p��莄LK�9�L}���W��$X�,�a�?����2�<�Γ*��+p_��N�1��x��;'�/�W��RZ柂W}���A�I?�ɳ��?�,�s��y���˷�K���?I���"������������<�����7�=��:G�R���H��C����ёܻ���_��������]E����n>�◯�?�G�Jo�Χ��#�w�/��@^@]5G&
[[�%w�ߍ���G��	�5�L��� ���nX�f6sog?�,�J�۴l��rtt4������	��m	k'�̗WVg����Z9��ι.3��5�P����/UuW{�Տ�0E����p%�5f��7uҭ��:�ٱg ���J,)�s 	��I�]\\Q����/�;�v�zq����իwiuy�3���mB�Ǆ[��� BLAP��&��$q�u�r3a��*�NK�	Ѹ)nn ��iei;mm����B� ��`�X&�(|��.������`�˿����Oҳ��t�ӣ˴���^~�*-/.�#��X"� �x
�iW:�@M�f�,�K����][����W�+m�*���J�4^f�!wt4z���{�itxXL�[pH�����A�C4J�P֫ʥa�$ 1��B��0���P�LV�̮�?����?�^|7c�#�*;=r,�p[hǽ<D3�Q12j���pL���Mc�nYP''�n$8q�!��luy��Ä���ݍ�Gڂ���x�aI���Q��=²��;����l�pr�brC�uo�;Z�ZvG�r*������M��U:<8w��ͩ�h`�n[\f�)w�:q�[V=��3 tNY���<�@ddt@B��-^�� Z@��^��x �[|�>m�ݴ��Il76����Fz�b1��s��j	�
^=�����)��D�e�)���+���`�g��!��D�E���t��{��a3��*=���t��9·GW����>��I�k�j�ikkS��뎊3�)�A��cx��|���_��̀��83)&bp�P�"���x�s���%��v���V���x�H�ru%��N\�<<�F��۠0ثg[ROO���z���x���f�y��������7�ͦo�}��ugw�y	�D��FT�����O'D�\�����|Uԇb�=�d��SA.���n.�t�.��YW�fq\"9��­x+�aC%A��������=������d60z��H�y�p�7�x(�-���0�����>w���������nC��Yb�7&p(�NU�7Q������lX09"ag3��]�G�g�k+8`TU���[�C=��UfE�꟏�.$�K�9��p�T{�8Jp#5�,D�#��_�pF��Zϻ�g�qb�w���Jq%����IG�׻���[VI�۟��y���{����I���ƗV����������_�&mo���h�Lp �:�6�!�8�YB&+�#x<tʄ����$xޗp��~���?z��<��珞/��/-��2�~=g�ywD{}C�n��?�K�eE��n�$��p;-�v|d �������z%��T̄ �omu]�ԼW���;�A�|�0m�U���e�5F��{`�C��CӪ�Z�y�������\oQ<�v7��#@_�ØP��:��`j��N��ml�K�E���S�{�R���,W��гeґ�}������~��{������jhT�F�Pfᘊ��%�� ����5��5�����GwUSi:����at,�##��<��1�ay���'��1��wr�i�~������0�lƧg*���,!�6�Nt~���*vc[4"�f+	�/�{�fgf�!����^O	1C��O��p(��T�,���g2$t���a,0��zXBnT��[O�F���>���c���otfѫ����QH��$��6��2�K���a�P�-$�z���*��9Ns� ��m����{f1�	@x�HX��M�\��Y$
^-8@��P����A劣�P�����$���sje���,Щ0QL�4	G��N��^tˀ�rz&����,83;z�:mO����Cu����ӄh��=������ �lK��=���Ă���s��&����<�=8p�cDu�-6�c|A��m�̓� @��0w��D�/8'ĸF���Q,x�(l����
͠G���j 3�v1PNǰ�}��Sp>�1�EaG�V�����Ĺ��u�at���
�(��a������}��"�է�ڲ�8f�C�Κ��A���vZYYJKK��.�.�u;2��j�w9��Uq<��`�r>�����	�/�-�We����?�J�O�O��������/i��#�p��۱�[]xMV�\^Іix�ұ�	���+����fZo�[\K�+VqcI�\��W��p����Pq���Q��t_fE�@d@}[w-�� S�����D��?P()�x�G5H�E���'ӣ��X&���������0�m���C�g<�ay���A	ƥ=�Ze�8>><I�wQ�w ��4�-���:�\���G��.����p��D-���S;�<���/8%��0u�;>[ر����^�l�a�!&T����Af�U&�$&���[uPmγ��2ia!��_}V|uѯ�u�=aTP\s�u�&���9Ǉo��tv�#��CՌjǪ ������ϧ���7��ɋ�P��_,��j��m���?��B�g�r�&&�D'�V���Q��DTuVV�$x-��͝PK��FVc�(0�}��kPEĞ���6��ϙL�Ī<��T%�EޗSԳh���UZb%Vߔͷ���sv^m���L}���r�$^����K�S`�=�vq�$����ƽN;dB��j�����ġ�?�<���%�����`��Sm	+
ʏ��\��_[;��������W�{iA���3йe)����[f㘅dČ�7ǘ�	�jlmjl��?{�0=}x/�Wc�U�21�? ������Q���A4̪u�.������ҾF .�Z(v�	R�ʝ�P{ .�"fQ�GO�fL�A�%�ӓ�������滴�����я��G��H�E<�,Kh�D-��(�;2<��4��G�f�푧L	]��X�PZ#���g�*a��I�XKSy �kr|\�q(�
G-"Zh����fz~H#��9�nscS����_t�0�ĒK�[l޿_W���QN�.,�2�\�2����6u������t6/�Y(�Č�i�WA���U&�HK-.t��Q���z�.��P�`@�im�ɖ�[� (�2P���ӵ>�2dTS~�F�mi�R=�j�� =~x7M�����=Kw�9��l��'l�C���(��>�8��Z�����>v��Ӧ���ht7��cBu��=��[6� #K��<U؅ʤg_�� �̯:a���<��زxY�G����ɳ	�eI[���b�C�6���N\5���pQ��8B˟���ͯ����Ϫ��LF&���g<t��&���yw��i��a�b����i��V9�acU���g�� ]��G>"dg�G����V�����œ����!�r%-���<?�q��)�����_���۾ޕ'� �z�}��x���3�#�i�|^^u����ih0����w���W�ūW�����̻������������c2 �8�y�N�Y!0`�7��`�U?�j��z������/x�����0���x�!qT^O�5V ��ܑ�ן���Ual�q@�VW�\���w�+�z��i��3�፨�g�ފר�0��YB��ٳ� ��b���|v,}G�v����e~�:@���ݕ�=9(��>��O��Ѻ��k���np����l����{�5Ю� d}`��o�۸������|��ٳ�@���8R�>�W�eA+���)j[�g~U��U�+/B��Q/�}~G:~_�Px�����6��>�q	�ذ��-��zcx�C�ӏ�����0��O�~"�N��z_Ϭ�bJ��}y���c3�񣇺���{`ܕG��������o�\���_Y�]^�L��-x@�ē�Hm��F�O.�iZy�3Q֣�c�t��A�@���`�M?�^=��B3���0`,,"��"�䖶V��Uo}�i�s	�rUWn+��H�ޓ��z�;���':A��U?�[�ڇ��H�<P���e��#��q,^�`�+O�:%������ށ��ޥ�sjٵ�ҩ'g�?��鐙����/�۲F޻jp��,ѱ�`�p[#J@2!����/�ՠ=J�;5��?���MOH��P�j�Q0�b�/,8`J���"��y�w[�6��H��r��,�		|�<}�g̚����dG9f��"܊�n��	^[YO�_����k��)_���	�|��9�0K
��,5b[S0;#p�j��0���*L��Xfha��fv�Չ�3w�n$���b�� Z��Q**�ٸA	����>�_{)��	cc#b�]�ԓ�az?��VV$�n�pk�Z|v�!+[�{�,�P^���/u�W?�GpI��iH�͹I��!�� �:���3�Hwr�#�Q	|�c���^L�Yf(�`s&�f�Љ
�1MhB�?����->ytO����F�0{�@��3�G��Ϻ��2�坘أļ���&yg��QfG=��knn	�1����A3���ιG�eG5;��L;[ՙt��P�>1��Շ��t��T^n[0&$c97TAq���â3�M���2����K �S:Q�a�3�r��`:�;:��F�_�Ǟ�H�f��_#؄PG����3��"���h�čg�ӑӡ�!ԲB�h�c1c�:��C��Д�d FR`��.�*o7~�!���ᤓ?���g����|����Aqn��o��������=�����\웎@�����G��3u��!z�lH9f�^��̀q���Gyѝ���)!	x.]���X�g�V	�b�e�h��~�7�*���] ����Ʌ1����p�SYa9;9Tq�%�6������O=3���=��.ŧ�U8���c����A�Y��HY�fB���)ɵ�M9ۜ���ت��_�G���(b�Js�����~��:�W��*���8�r/��9Qތ Ǿ���Ƴ�]<��K�kk�ikc�3��nQ@}�W�D���L3\��p?�	|��G�l$4@_���y�;���{��%]���z��'Oŷlr�I&�Gf��Sn�����P�c�vlt��f�ś�z�۞�<�:6�A����v��w�k;�>Ga,�3�H?�LE߼�����/y��2&����TQW��f �L1,f�nY]�0��`H���U&ʞ����m�+�  G53YĊ�y�wnE���N��F��1�"�Ȯ]��-�ˀ���o��|/X��� V�9��G8㠬����B�������:|���_��>�+p�l����0��bai9mjPv�o����_|��s�VW�d*�Ct���Q�N��p�и�`N�A��;91��2�PA:������f;�k��i���mW������ԐvT�iyi]j'� ��*�,c�o�@� [�̴�)��:�w�C�eJ�ΟY,:�����p�'|=��%���7L	��ޱ;6��eٺO�.��V�e���mE�p�Fl\b'{��" ���1�Hl§�MHpt�2k�F��'&$�c
�Q�r��b`I�f#�C�UV]jtxd��e	�±�X�P�q�ĸ#�p�^&<���DmƢ ?Ԣ��Y��{��QZ^6���l����+M�~j��������c�{����2*����3��e��Z#�X�����1�_fK1���8�o�����M��@`~n�;V�Ÿ�v�=��Q�����N;ۛisCt�g�w��n���-;ag���lthe���x�Xf��-H�E�Y�N��v��q�)I P綻��vՐ���w=�*6��\���F��\T�B�G��yg�X��R;�V�)�T<6J"й]M��&�FT�Ww�h7�L��>:2g��(���p��rB��otp<E{��s0}ȉ�
�}���j�WҢ���B�������u-<����,�����~�o������ή�j�)C��O\��^/�?�l����.3�!�b���;� P3gul"������������-��T��-_�� �J�Z|ɳ�tЮ��a�噭ҵ�I\v˗|LO��l
���}��y���!���3�� ���=�������V��"�1�knc���7&�P�`7�wի���aĞ�������~h]��2�"�q"f��^�!5��X!D�RV��_�ٽV��v��O�(�.���c	�D.�7���CT"�K��]�n� �;�$���JZ]^�ҷ��U�M�klW���!@���k� 4B�*9�����g��-�4��ݑp�	�ucQM�U��i��~��ZD�6�(�$��'��0b�U��6�We�7L`>��tQ9������n��noXB؊p<qb�UF���?���E��n,���g�'�#N9�Z��NZ\\mZ�����?VnisL�1��M���^O���Ȥ3�g���f�1B����m�{�b� +����E��� FQe@�a֝xVq��Ʒҋ:ԕ�˾�e��x��z�T|�j�xXتe�w���ԫ��zA�?T��V�-F{+�o�hQ�u�����^Z]�H��˶`�$X��o����e�z�W�����
�"���	��%lR��/�vԺ�T>�om�Wogӻ�����*�k�B׺���u	`�2ø.�+�M�1�ExaB~�E�֥�ظ��J��bC����UG8 ������@�&0BaFtrjL��]>�	.0	DF#AG�F��!��a�f�Kuި�/,�
�b���@��;��6��Qi�9bp9DTg�������^.�0��c64�� (����AH������4���V�@�G3w!��HyB ���K�=qpՍ�Η�HT_�������Pd�=������ٻ^�ᙑ5�1�sd�eB�K̢���=�h��8BT�R�{:��{��qt�P���X
��E�{�j�.��'�"��a*,�q���ގ�m�������^6�F=�K�fh�f�#���:`!V¬�%̲Ⴡ�y��f���۽�ɦ��� ��Z���m>P8 �7���I� ^�2I���J�n@�ε�_�Zu5Ѧ]W��̄��H��ÊǙN�}���tp����!be��:�'m�A��+�̘pD53$tX��To`��l�d����4Óny�k�:(t>%��\��r��gp��?WR�8乔"�"�V.G�w��=�Z�
��c?vn�%�޽w�~jz:�ONY������ޑ�t"�#aL��f��U�}��$4�:�)�ϯ�ĩ:��|��'�"s�r�p�֝m���=g��`Oe��m����� ��%�nq���Ev��~�]��tȦ_��M&4�p� :L<��#�9�C 09u�>f�X�\�3�/U=�Vx$�X�t�L�">ˀ�D<�@e�`yo_}��]	���bR�~����qlिb��Q����T��2f��ݷ���Y��^�'�ߡ� Ϟ���wx�xa��H�V��Fx�X),�J��TƬ�p�*q�@ވ:�a
��{�e�}�|_ڔh�X�!����x��?a_����F�܇²UY���l��<����+�w��TA���M{�ND�o���O S\I�:R}�%N([Z\W���T�(��H&hP=�d�Vh�&�j0?{+�]�?�p���YH^o�-���@�W��C�?)�A�eY�� ��{�9�1V��/s��:*��<�:q�%�k���z���������j�`��0��$�K�vVx�����.�U������d���5����F������H��Lvm�S�q�����L$�Ɇ�1��V	'�1#)�AizN��_�}z��mz/f��>Ć����*�eF�\�"���-:#������@�ƌ��!(,765ņ"�,1�555�F%��+˒?�Uf�VW�U�W��Ť���Ԉ '���s�ŶG��b,}6�@Dhj�T�C����I���&b���6�G0Q�l��X`>�@ �^i��"��gfU$`�"�1�͆2���
G/����:ck�Pƈ�G�ۍ�����|��-�<3�,A��cPƨ5P��𙱘���� f��߸��ы�w|o�Q������1���&ӓ��S��w���`��^F��uz�@ �g�WMb��O+#c��4�W�/�)�)�	m���-4�	G�X��;��o_��%4��7zσ�ARv���=]5�:A���	Z*/e�t�a���5gc3�����Ϭ1j�K��f?��� �)�,����J�+��Ҏ�%t�`2�eD��05�4b�b$�t! ������[����C,�-��(R����5�c��}"�G]y�=����B	�!�X�,��a�tL��LOMX݄����+�� �h7D`��-���������A���[��N�n�����H�/�U���ֹ��(���êļ&�/����095�>|��=�<=~�$ݻ�@��4>!�g ]^��Vա�p���1�9=�I<˫o��jyyڤc��cv��X ��M�j��nU��R�9�:�R��o��sa�Vt��X�~������"��N�{'^]|��eZ����Ѧr0�����c}emM�yC�y�t	�a>�$lmu5mk }���@��?�^'�	_���,�7���G=[��P��K+��g�G\w����Ӯ�'ƕ7xE�a�̌�����[6\3���y.��I��o�|R:��w^�J�l�sll-��R���%�Ľ¢�}�L��wзeeE���KV=�Y��M���O�ˠOU�M@������� c3���@���1��)���S�����??8O��g����y��R�B���ӽ�(������Pur�>Ltt��l����?��Īꆅ�s�qt����,ܪ�+�V8Gf@^Aձ^��Ĭ��rۊj��D� �,�YX���&Xpb���@��P��&�h�M�
.D@����o��8(3\���[�g>��`�ʤ��<;�ח�U���.�(��m�K&e�3�����"�	�\+�{ie�Y��4���v��/����_A�,�bĘN-�"!5�!�X��ñCi=J5@f��M��%	� } arqy-}�ݫ433�w��{�As�8a7�)	G�Rp����B0��H2jAfFv�/�[�WcB��͘IA_�P�7���6$LS[��2�76�j@�F}0���a�\B�D�d��� X�|��!�Bb�l���УD}�� ��`;�K	D�~ς-ԩF!e��C�RـS��U��]���u���Y�=L�e�^�e$	�ʻ����3u�0��5�xt��.>���r��ZB�E�����>~|7=z8e:��$�����G탎��Qݔ�>�L�[ԓ��P��N�8�Uk��(�3�a�F�q��K���d�!3��Oed�p��s�j&�V!�B��`B��4&�X"bv�/,[�A�����`˽UZ$Т����f}Y�U�Xa`�����ع�`
�#::�1'�S�l�������=N���3��!P���{�%	��RWٻ҈�]�<�\���X�p+^�>򽃀>/��w��u��`��##�@���)�3+G�[[iof��Cu��\6�4���$�p��#��H�q������� �TU����At*QN��M���T%.qHC�.L��x0=2:&g*M�c�̤M��%:Lw��;Y�=Jkk�8�&��X�5
��X����8�&3������(�lZ���M����y�ªw*+�N�w��g֏	T�P%c����>�J���_��d�YJ��6�S	�,��{ ʄ	�%fQ]`b��AV�X�A� '��#!���G��<�n��-<���;�[���\YlR�Ky	C�G�ܪ?�����G b��� #`�!���8�+	��n�k����6�bZ�{Xxy0��̨� a�ዶ���wb�3�#�؛b�s�����$��͚��@��N��ć�e���T�M�6*/�Wt�{��Zv`�Vx�����#��	���X�1������J�ʿ*����U�?��P{��U�Z�sx���3�n�:��kT��'��N��mT�2����K��`
Շ���eb��&:��E�ܰT�L�)J(���~o��
O-��!�2p��^V/�-��E=���͎��IQ��J�w�l�%�\�8Ѥh�g0�����w�&����ْA!'�^�|Cé�w ��N��������;�VIX������1�����_1�d��@���fF �~�g ��E�K �8Y�M�"l�ñ���ٗ�gT�k`��4?�n�ތ`��L ^�lN'o�L��U!J@���2aˡ��p�0n,ܲ�?�f��Uz���j�.�-���>� �\�}�8���l+���:�ª��%��U	�Eo����X�D�`�	B2�dɆ�t{��#=NAf	�S1�c�ak�����j1̭�� �Dg�Z�K�]��ۚpˬ���*�����*c�ӣj$�h��z�� �*��I��B����衲[�lO��K�S��g��iZXXKo^ͦ���>}�������4?����G�+��%�1�,.�Z�mW��Ҡ�|��~_�752�����
jt3�}�(:?Q�b��pz�p\�R�e�=C�0F�X��̈́�R�#�S�Xr�c�	Y�@�+,B-¬���=���m�\\5j.��0��(�&l�12"ZIC��J�%�wR0�hXH`Wt�����s�i��M1ޢs]	�ԏh�&DV(����#q���\����x�."�_�f��N� uN��)FhSJMn'�bjX�X_�߰ps�qC��ô}ճ�Yde�ƽ~]�Я�(:����?����#UP���"�fO��}n�7\~,�����%:<;��=�W<i`h�˄��/t����Z��,Kx;�� �A�8V�,x���b�����߀���p�ǅ��_�\�ƻ�w�'M���
BC������-���9��_No^���jI��LN�'�y�f�I�젣��ŝV�C��i� 'Z��Q���$}���Xv6�2��5��#���YVt\U'�0X�a���4iK8�4-f�8|����B
'�݆����vw�.&���#lt�X�y����5�~���=��iz��az�tZB�xl��,��X>����8jw�*��
���N}#�`���&�;t���;��
��^Te�Ъ.�ſ���G�ER�!/�A��2V�N<������Z�?�fgߧ����{�X0x��{l�����ev����y>޽�S��4��i~��c�W�����33�қ�3�;�gl�.�Vl�xyë�#�P�;�X�#�_��"0�BOu6V��3������؃��(&T9,�XT$h�L� ����>�3&op�:�$+�V��n��(	��KdE	��	�Rx�Av�x.�+���,4���L��[�>=��7��\[fݻ�������^����**��ĺ#�nU����p��%3�,�ȃn��f�s �� =S+l3ڤr�8��+g!#�*y1<M ��+6P-o��u�����IFX���t�8©�2+���{{��PL5�;���tr0Z/�^/�#,�	��T�q<��=a�	#��CF��^��g/ ���� �NZܫ��_��+@�.����_�tkb�x�j�u9�>W�}ݳ��+��k��wt��h��=�����=�G�d�����b6��Wߦ_�����_c��_�&��Wߤ�mF��:��Nf�8�f4���]^�?�8�H���� JW޵�	tvh�Ȓ����<���@�λn1e̴!�"؆�Y6"��[�q���i�`�S���a7A;�y�j]튇��H@Fk��� �A}h)�	aZ4z�9TS�X�,>:����Neүq��+\>j>���"G��Ϯ���+iW�8���A��\}�gys��@od�+7v�!Ȳٕ}���p���ߤ/ި#��@g�˧��@��Tu��M�=᎓=03��W8��%v�|鷻�������9Cl$f���|k��'��+�_����G�����G��#�HK踭'N�\^ٖ0�}�#uR`�<U�̈2!B�ƕP/��sA�$�?w�l�}�������l�t�V�0_�}������9�x*!��V�� Mw�x�7&!�@]2ISh�#�! #X�_�0���lE'��-��6����vw4�>�Aȇ�屽�I��v�6}�A���3|�:BsÕ�)u�7i��aw@�g�u �3��4{xǷ�a>��yЕ�{h��D?|�8a���{0-�MX[@��  ~��B9�w��	e/N��~V/��rMu0�s�J��}m7��x�X���ok�
��A?�����33��ի7��׾�� ^����W�P�|��]z����������+�����{����^��3�C3��U������o_�����˗�%�Ϊ}�Z]�v��M�1��)��(��.�X�C�<H@w{{/mi ��/A�8V�D̩Ai��S�1��YR�eL�����W��Ӳ�u	���W�++��g�\�m��a���,��_�_�Tp���HxV�bb.O䴉#���a�tgg��JؘIvv1�ۛZѳm�$�PGՏs���{�vW�j�/ԽH���=��ka�2 �Z�����\UL&V�56K��;eR8V�q4kĉ�*'�1���n<3�hV��'#�"�a�<�$�c:��� d|0��˳P�u�NɅ��<*QXNM���� A���A7�:g�3n1N�P��$��1R^�G�QO��4!�f*����<��yiը��A�]���F �Qt�Msrt�8b��M���6� $�l
ϼ+�9�N.ڏ|u��ە�*a�BQ�۾��z,�c]"�3ԁ�h�N�Z��Fjq-.�9����̥���4����1�Wb>o�Z���;R:�0M��f�:��Rg���ș��Ij��5"&�����:�]j0}b��u]��)[�h��M�ЮN ��XX�CM ;�����,0��3���/��mܫ��������q*�,˰3�Y���9b9�Q,� �Z��L��~=�!/Ы��C[�xѧ��kd��:�W�!	xD,>;nK�W�^����},��]N'R� ��}_��v���鈴�4�tؼ� ��_�*�������?N�������?K�~�"-/�$��{��Ҫ���oz�����f6B��Ź�`�;.����S����m���S�[�'���^��z��<�����v����o��o�K?�ٯ�?�����e���ߪS�W�]���3ڀ�������٥��� ��U���Sg�A.f����3�ޏy�r�Л=����U���/�׸����:�{t�ᳬry����v�Ҧ����C:��6��r�Վ~�.��&�&���E�T8��b&����=�!�`[����됄ٱa	���i��O��5��0hչ�8(b�O��K�" @�����g�{�����nyf@YznS����YZ��pÓ���O4�K�����M�spʊ�� �ot�Y�;�@����^��M/_ͩ=n��}6�]i@��?�y;5�G֠O���Ө�uzьjP�fϽ�8O�ן���
�q;$ ��0�I)VZ)�P9��
���+�&��!�P���0+��#]_ٔ�J��ljB��B�*9=�]���-�����t�����xE	S���������cV��_L�*3p�<�5��k�΢�V�p�}������%ViQ��ܱ5THH\by����P�y�D�����1S:?���I🟛7���HGt�p�~���r�z,���'���g������P�~��@�Ì-���觩0Ll���lY�Œ�!��ҾгU_`���jˁd���]Mn��T��(OdAHg /���5����sA��� �����:+B��*�)R�<eH�e�D�Bm\��~B����oh]��7 �/�σ��AD�DD/ǣ���X�gY��0v�<Vl8ը��Q��X~�Q|�g",�Cy��h���x�z{`!]f��.®����g�	7^�K��;1�q�x��?� bC@4�}NȂ#QH{�P��O#/3�E��̳Q�?2��z��� �/ *7x�Gʈ.�����}j���b� �!����UD��P�r�:ł\^�t%.��J���pL���R���y��m�pۭFCC�0TQ�QV$6b1�4�0�z ��E�3L�!	�6�'���k���Wˠ�ϝ��rGJ[�3� Z7�Ԗ����PrU+��e;L����4�Ͽq[����e��L���8���zW�ׅ����\�e N�G^�KE��R�qt 9ҘA��lz�� �����ŋ����4���/K�o/q�@�g|O[垶e�,Hr@���+�|�s�9$�[�-^�����a����q/W�U����C�%����իo����W�7_�I_�L֜�I�U'� G�^i��޲
������ȗ�����"��GT�u��x�ǼW����G>p�;_���ݼ7"�_O�(,��l��Ft_������2jc�[=����+E��ӻ�=��2��%,0i���|��.�_�q�Y�t����'A�Y�NyV~|�Ѣ�$,H@d��L˝�I��70���6��G�+w8����A����2��
���b�}7���޳���@�2#Ľ�y�~���xՍ��U�zO�;61���%�Y�U�s���a�+�E�C��"�LY�Z�^��w��tI34���U0�i����X�AEp`H�
#-Ӛp�k̅1{���m
ǺM�uV�j�`u2�tҿ���#<(&��� ���tU��rx��pU��@+�oɓY[�z�Wn%�o �G2�`���M�*�Sy��P�B��Y\�S�a�4�%�����,'�"+yfX3����&%xm�X�c�O9#�=��U'<h0��Dl�֕A�jC����ؼ
���������6QEРK< �3�[d�}�.�~�jʳr��^���W�l��o��,�2dE��3�z��,��ߩZ^^�B�۲�hA�$a͛�D�(�[����a&�+j�`D�7�ʾ���s@�W4�\@4�a�Lck���mGR���s5���h��$4cI
d1s��mL�C\|c�2��=qt\�QB����9��w�֪ۀ4! ��0�B�����I�!��p�.��\^�kt���VVT��ra>ԑ� TVF=x7�<�FNn�bz�q�5�G�������C�)b�ȡ.��Ax�U�C�̌E��۰l���Ck4��,
�����4�k_�������t���t�ޣ46>)ƃ��J��:�C�eh��ިo�Lpl�
`�UVF�lТa[�U�G>��7ywh��l�@��*�N6e��o��:� � o[��j�!�ƬR���+'��tͰL��]j��T3��;~=��3�.�/a�Ұ������4\���W�!�$�����J���gÔ��G�c#W�8�:��}��Atv2=�Խ���{3"�3̲�z�1��z�$�t�,cs�����?�"���Q�t.��A��>�?.쪭���HA):?��מ�8�Fq�"�en�e�����l,�J؝���[�=�p� �c���o�!�*�,\��(�s��.h�#!���}~_7फ़�LU*�g�<�,>�<�-80n�͔M���:I7f�\`��X��N�� =�K���' �*�f����qB��*!D�A����CWN@k�0� W���󒜎�;�Z���p�vaa�'8�E�#>gЬ���Ă�y����2a����q�����۷������ia~�3�n_ʏ�	��|�m��?������闿�ez����}���R5T�:r{������.*����0���I^G{�O�����{^T��Sa����Dz��A��G��O~�E���}�~"���#�'�����JC#�H�Hqyw��]���w�o�A��F��ɓ���8���A��?����)߽wW�ِ�n��'ʂP�_X+�TZ��u�~�}��y�>-L_!���Զ�v��p&��%��JB�gL=`���G���y��l�J��1����r�f��`�/xc��k��A/z����mQ8��1�K=#�	��Ɋ(���]�}�����+�CC�p�v"��1�=� �Ѻl [X\I�痬#͆�]�����m3$�2�4��B!�XFJ�+�+3*�d�lY��� <]~p�L�ln�J� ��d������!f,Z��g`�GWF�00�D#�P�F��7�\�����e&0�n�[	Y�Pp2ˌ��&.��I�el�g��(vwb��������	<����҃�^�У���������� �Z�U\�8��aw-#sODy�@@x°9�.v�7zǻF�b�[�qY����,S=nuEu^Ag�Y
5 �Z��W����@j���n�d���[��v����C�n��NX�9=��ì��7�%V+0���G{��g��d��+B5`�|{�(ml�@���|<�ѿ�L H�-�I�D*�;r�Q���*=EG0}��X�D`�t�>��8���i�����^x�@)oA+_}���S:���Y��R�0�`��;�0��p�"�\��o<;�zW�av�����]}Nd�(_�7��/?�"���х�˳���D�e�I[&��f��k�s%d�
|�ĥ���ԙ��r�?��~�����s$\=��E;�����;_#"�3������z�
�X��mna-����dW6l�q�M3�o��,O�GYۘ-Tj��v,�4��eF�����RW&�z���8p+B.>�n�]�b���(e�WQ�ޙ�ĕ�p��N��;��Б�`_|�4��c�<����S��JӀXP��)*Q��	G�c��J0�Ƒ���p���k�F�'=&� @"�"� �`�MG�	 �5rc<'!���2�11}�1n���|3��Q�h�k[�<B��>pn��
ߊ��gQ���x�m}x�U��Ņ^@}%�-����)��wjz,=z|/=}�0}����ŗ���O�Y��G�$�����~	�l�Jh���� ={v_���"6S�ꯚ����?{�~�����/���#4��G��'O���Io���(wE�*�W����ʀw��+u�0aJߢo��&Vɱڰ��D�.yk���79�(&�H+9�\�H@�)QTe����P�LHQ�`6�~���Oy�aƘ<`=�aj��yǤO��ec�'>��f�<�ʘ����� �z�#���0aU�C��QedS��p]tnOX��� �>D�*���q���MPB�D��_*���;}�Ɗ.>�U/��]�	1�9�����v� �'������V��wA�sV�i׮P������`)�:.w" ��Y��t8��G �;1������lgJc�����G�I�z/B��X]f��%����C@�%/�`tf��tUY+�l�X���=TTn�^�����aW�o��{;ic�)��
D��jTU��{pF' 13A�W��7H�f> d  ��IDAT���W�n����>@�n���_@0�`��s
jTf�4J1ofYa�]���ޮFէ�ws��5�>u mb�l�8ݴ%�f����a��*��[���."�Qz��;g僐��C��2���� ���c*Gx��1�Ƭ{�vK(���Dg��a�d���8�g���^�=��Yr�:A�Y}�h��?=������3��*K<*o��vf:6j�'��9�rt���x��E�.l���?"����>����#��2>� `������끵�h�L)���RaW����������cpn˽@r�O�x1nx�� %�����.������x�e�z���@�W����#� �)X^I�0�����3C����K�j�	���ō~�5JM+�e�6��C����0e�vۓ� ,@ӿ�[��Pw�>�-�_<h��\p�d�Zb
!xH�D�R<Vcbf0Vg<���O��B_�cT�ˁ��"�2�{*^��3������?:�Q.����!�
9�h2\��޻�[ZR��6ĲO�w���蟙)��bU�}&}��!���%p/���^	s�idx$�Ѷ��n�׬6ۢ~���2#ihp,�{�+6���E�UVP�ڢ�[ �y�].V���T�<A��݊�t �-(��)f���G�m�����?J�}.�Gӗ_>J��{O�O�H�|�N��O�ӳ�~�/�x�>{~7ݗ�;0��:�Nb%�9M�+�Gӊ���,}����񏟧K���ϕ�#�YH�!�M��D�u�l�M4���2=@�����(����1Xž2�T�£jW�G�$]��	K<�lfF���$��f�a�f?m#4oq�.�b7�W�j�����{S�g����Iͻ=Z�E�UT�:��8�A ' ��v�]��BM��h߽��f��܂d2ّ`����tE˲j�4B�+��(VD3y����6���Q�&T��|���a:�F#gS��ɡԱC�y([�H������miX>���vԏ���j�p��T�)b��ϔ��0z`׮LIP�&�,ַ��@PeW�MM,K�P���h���t���l,��Z���L85面��<���{�f4���_��6����e�Y����[�'�Ęx�ŎB�1��b���J���*����p!xi�\jn]J�Y��T�oo?;�8 ������ �޾�p���M�aG����51Y�Q���β<�,q��p�q�^���jz?��ε��F�M��4�6P@�e��FD�3#��]�����&lA��'�p�]�j-��s-.C��h�yҀ��c��u*B�p^N��+���mXD#ć KY�W�KJ0��?�*�tΥ�sU駾�/>^��Qڒ^ ���A������:�ԢU�z�.�[�ɳ|j��Y�>Ӛz{���g����Q�Ruw�`��c
 ��W_�sx�[�g�}�9,��(o��򸏅g�	����W����ދ�~�w�+��k��\�'�N�����٠�z�[�Ju��yB�2m*��E#J��'��z/z���-_�q��E7|�K��D������"�W���O�e������[_>����+q��� �%VL~�]����M3��>�V0��c0l�SN�>|���l�X��g-3Y�����~}�g�{�P�Ni�ɍ��%̺������:1���Tڦ%<��1=���N���1����Ơ���C���O��/�L��}	����K>��9<BU���������"�h��S<�T�r��Q�fP�s��i_�#LOO�G驪��z�0&95H���uh�WeR1i:���ʏ��w��h����p��a��S�a�-F`k>�Hc��<8���N��m{�S���O��A��=Q�q�U��>r�vO��>c �f8���uy�B#�b֕Y\��H(d2-�/�2���\��(��Z��+p���*���q�'L�1iy����i��fo���J��5�w��BS�)��f��	B�xfk[�x�D�B�Zd������+3���k��j�}�����7������J��w'����@�x��Ԧ��4I��KO�<֨��d>Kϟ>N���\��0g�zr��Ύ�q'!�KD3���D�gjE`��GG0 NH�W�Ùa�E�7Y(@�K�uD5�X�T�g8۠GG���I��� ��
�Va{�'is{_�,ǻa�e�mo�Cυ�*�]w~Ό���hjm��������:��gz<>���{�8[i~qE#��43���%Uؖ+��u��*B�u{���C5�����R҉G�!�Y���ڦIx�M�@�Е�kz�	������H�=? ��&<�fa~-��l?3�W�w,���]J��&}�����y��cq�� �+��Iakj��3��o_�_�����_�L����V������`��=��J'���Lx�����p��ζ/'�r�lR���h(�J߃%<偾�єN�q:��Ysն���1��9a�p�!}e,H�Ȕ+0�Ј�Tq��răU�6(<������g�E߅@�N�:���!�J�R�v\� ��8�+����$�����~\V�`��Y%E(�ƅi����t����H<���ibj\@���\�9��q�x�JW���)O��3wdĿ�����V��b�)��k�<��>�ۤ�o��x�(C�wyT��N�Uނ�-_�em�4{��\��j�`Ѩ��j6jm�z}��q�}�	&v����I��6���=4��ÿE���G�wi�F}��'MeAa��,�E��Y���Eu�5����5�AE��?j!6P�hp�����������?�h�Mjf�:Վ��'�tzOYK��>��8��&����ݽ�6`��}^�=�{3T��L%g�J�c����e��+q�,��8i�]���l!B>T�\@�9tt�|�G���ӳ�b�}|j,5+���&5K@���>��'���_H������&��=Is�z����g�W/Y���|e�3��P�r�7�y�K���;��v��7/*=ʉ}�)�{����41>,a���� =U�?��3Sɠ�&%�K�E�%��e�Q��D����p��F��է�" ���*��p��8�mxxH���h X�",��4sJ�Ht��p� ��St���]䱧�l}cÖ,���_{��e"���p�j����8�����A��ب`�``�x�^ �/���������{MP9�� �9�'��x�M8�0�|��O�<8ȁVz�O�j3��Pea������m	�Q�%�`<�Bľ�It������w�M���T�4��Tj̍��#Ct��Q�Bե˨FCS6g��gz�#������`��jO��b��q �t||0MM����Ǉ�mD�!���]��+��y���L�����s�v39�D��9�U��ѣb�O�N�	�R��v�X��6v%�#��	��l<��|v-A
��BU�������A�6i�s�8M�O��7��M�T���A�U��ʗ�7��}����F,\���1���\v<usS�i�NΝ�@E��jM����"�q�WPW��*��ĳG�e��US�
��������d���	ߛ������ul<��9�3'1��$N�F�gj(����w��7�y�^|3�fWČ ]I>�V'�46:�hD�k�\0d0C@�Ű7�{芲AA���w,�����(����Eܳ�A��I)���&����<B�X1�F]���L��X�3Ƣ�MGo�uh�q��C7���ci�u/��#W���������L��
b����	On�`B?�.WyUw�\�p��ވ��۫��<��>�&<d�8��E��?��N��:�i�u��!EV9N$Ȝ��"�^�G�-��*�7�1#[t�G����l0�2;�o~���x���Q�zEPx��tF|J��4YS: �AZ�3ӽ�{�̕g��rx���st��8�����H�c{����%K;��u%�vD���J�:&jм~�.�W������a�ޥ^�",p����3S�G��^iZ�5��{�������{��+�*g�t��~�N����/|��X�j��H�3MA#��@u� 9fnQGC�I��
槰���
�E����4.UyW��\�u ���0�n3�"�3�8N��*W6ӑ�x��Lt
���s���5���QB+�n $A�I����ID6�Q*��P-I�V݁'��I��?0����R���˴���f�V���ZZ��W�$DJ@�`�Ą��>�ms��9N�;��71�$�L����2�&s �e�<��{�0��®��
q�V@M���}��MJ�ClkoM�����^~�6}���ۯ_��o�=1u�����μqLB�����X��Eb~����z���/mQ��Ki�]][��N7�O= -<E��bx%��k�ó�P��e�1?�������a6D�r��E�S}�l6c2ni%&�$"��`\j�I�v{��V$�vkP�Ջ)56^w��d���@:B /��]�MK�z@5�U�)�'ZkU�=`����>�	'��_	���0qH�K晙[N��ӜM�m��^����=��J�n��8�0x�W�������b�qc���z1p�`f�3��:uà#ƚ"�+l�A_���n���ңSiD#�V�p����-����:t2�i\��w4�D��Ê� o�ihU��8�8mS��.����������l�O��]���N	���j���szz%vۆ�WVV}\'&3IQ��.���0��ʹ�{"l�I8�Z�F�d�z%�6�(�-�"��Э��!�ɕF ��i�.7�# 3��l,��t�2K�U������܂OUYX�W�gn��<36>&�S��FMz�"��-3��+3+M�?fl�4��h/�C3E����T�wo�pp�|� ҽ� ���%.l�3��:�=����H�n��qb?vt��G�Nk�î�K!{C��մ&{�pёa�Y�a�ȉn�j$M�Kz��AU:JݬC:Л~�~�34��� ��{�j`�܃��K�2p�
��pc13�hR(A��Yױ ���t�3�:B,�-�4Y%vs�O4K9�"X_���'�Yfg�(&ft	ds&'��J�0�\NC�m�ӝr��*vE�t��c�3�(���o)�B͠ 4Tn�S�Z��͉@⚽�<�"\�B��]���s9�>��3{�A�7�y���ܹP}u�{�9v"ML�
G-���s��zl�.YՀm��%��Pk�T�[�Y�F'pt: @u�@��;æ��3�LB$<��I����l���E�%}��w�c`��t~tR�{�k1$]�Ia��cǔ�^���4���%�k�Ku��w�s��Y1\�Q4��:{�QڗZ;��O�S�9,��_��# `Agx��h��N:$�l����32��f����谀�3B�C��=����Y"խ�f�O�+�%��~�8P���_�@G���Px��n�HO���q���B�w�(���x?;�vx*�iP~T�kDBS���d��8�8 a%�c��Z[��!:�]XH+�˝����-'Kr|/��� s,�,86�7�XV<[G��N}v���r�c�q�I�	�̖3��#!�tmVy� ͦf��Dϑ�3��������,x��%>21�= �R_�y��E	N�l�0HW�z	<���%�[Mog�=��P$����Q�+G����w�Q�D�sRyj=��8�	|��t�,�ڝ��x}O�wo�'��HN�<;M�$�~���������o^���<3��⣱�U4f[[;�_ww�&�!�a_�PX�a�sk#-.rz�l����O�F���cM`eeW���oyͫ�Lh��`="#������e��O���ojw���4*u�ۛ�O����Ѱ���@}J�z��J�]X�H&ژ\!O,4�m�L|�*�:��ᛱ)68�!<<9[�P]a�v���  !؂���q�Y�G͡��ó�xZN8l���E2"�9aL4�L�,Y8=nnɇ�����#�c�b��V80��R>mn���ڿ����:C�[:\�ΣN58#_��p|�	�/.Я8P!Ҩ�iu4$�b��gcS�u�b���C�mnityو�A ��9M[b`���p�zԃp�g?�WW�;:	����Tc�N����v*��o߾KK�Kj�k�F),�������]xl�b�U�$02�)��0����eY }v�� ,�	O��\܃��Cv"�c,P5@��Q��p��zYBua�]�W�Y[]Uz��א�<�$�L��Y���������E��0��鿓w�  F���A�ÙiPs�W���o�D������K|��d���=���p�9�"/1���鴅[L� 6L��B!��B]�e�k�<�ƔЛ;R�jD���@z�3�,�R4��Y.B���p�$�q��C�9ٰ��	�-:5�bm�D�����c�]�0�T��3q記��U��Æ2xT��cf�SbP�������0����m�Q(h����ޞ:Hu��L��|aR"=��q�[`�����Hh1w�=3;Q�t�J��r���&��3Q�ƪ.�������R!��w����z��M��@O�L��-a�ꘙ��{��c�<�Vu ��H��d�����,8��5O0���mk���a�"�@��̚�.�3�� ��(6���&�.�#��ol�m�wV�������E[:��4�:%�Y{ڊ����C�A`��ai����\#�>�[�z*}�>�i �,�ݛn��<m�PB���b��0	҅iy���Jg�w����a�������+zj�`��J�6�4��P١���wށy�a�(̫G*#}B�ԃg��M�:�8���w
Bǒ	T.�S�T)��� ��nML���h�p;����>`�;����G�=�;<",�vlLi	���C� l�b"pX���b�w�z��n���V	Qeb��ee��c�]��Y�Y��hx�?�J8�FnG��P�K����z�τ�@��=���r]�\��2C!w+�BŜ}>����^��E]lG0(/��z�`ac��{	�b����0��^��߲����Vœ���A�#���+A�#2-&�<���kO�� ���E�}��3�#$�F�.�}	��#i���j(�<����O��G`�V,xF /x/��3yD{�?X^�0/�`�]��c�.�{�%�s ��Ktw'��N{�Con�6�W$<�G0�a������l�okk�Y��INn�9F?��3�C���l�����0�J[���V���X2���]2���R��3�j9@�r�S|�W�?6I澗���*`���1���: �2c[=�_��1��L�/�?������
+���%�L���,�ӷ"؊���C���\�γd���o�ݯ��3�Ӧ�)x��3�VEԘ��L/�T�|����ςM�LxwB��QH���|���M�yF�B���9�n����Y�שEB�Q�Xg�#"���l̬��s1�
*F�g/�7�`�"��ӓ�'s�ْ��a���<'���{oޮ�W���H	�EʀeX"���s0P6`�{��'ib�O(��(A-C����U{����y�.3���W���s2�V�	1�Y_��+V�h7�gM�J�
e��>o���o��A�<�ɜ�ڤ��a�k�����x�ݻ��a���.\
B0ؐ��x�FK.�(*K��p�4y�ft�f�g�� z��1�um�hP�y���ty����o�E)�M��^8��o�_�v�׌2�����}E^%�fna �V �= !Pn�=7�hj�wf�Ʊ;���0�gǀ-S�$�SG�ͨ��v�W����,�ښ�D���.���%F�ڏ���>�y)�O��*5*����kޜ�3���GU���c(��䓏2z[��-���{����t�QPݼ�r{"e��)gҽ��1��.� �^��
��rF������x����fO�S����>���[`T9͝�T�|��z���;���*�j�����*�%�l���C�8?���b*�6�;ߛ�
j�n|�G�I
�aui��,���5����#JLw�o�;E������������ĻG��s��K�o����a�t�<�����~��)'�l�e�,u�y)��&����'��KcΌÙ�/f9�ܒ������s(%�=SA�A�'|l�W^��
��E��J���v�*�*��=��l��}����2@�����\�9u�tf�c�yݔa�Y����q0���
rg;�M����q	��w�viig��̜de�D�$���'V�����v��1y�2�
���GtW��Sg�L�x)��U���Q�"��%�NKYP_+Ȼ3@yF&���C�;{�5�)Tu�(2s�d�ae����:rF���G����7�z���IǕ��U����|��?i�$�q;s��/ϐ����^��r{�r�U�YZS��p�<*���8�V9t��2u��9}�Q�ޠ��p���|�z�[uTBW�&�״��U���}�w�ڟ���)�NR�u���"aN���3��(��ًQΜsy�tf~=t�ޔɥ���[']��Ǻ�t���鳧�d��Rɫ�"������Y�=��w�8�y7W���y �j���;뇾��N�T�^)��Y�<R��J���ֱ|Q<QzJ"�����уQn?��V��@د�9�n����W��.[�39�n�m� :Ab�p���x���A�z��g62�܆�UjO�O>�8g �߸�A�������w�-0<yN��� �UB�¢�
�»n����c~y=�28_�x�2����ۃ�{��*_�r޻��u�]A���u��Edׅ�{�-gEm[*��!��"�=��"��F��ֶςRlk�[
���2 Ȁ�̀]��6�U��Rp1�l�'m�V62;{�>��r떊�O� �u��J�(��O@����Lp�NǏ;(a0�����]�u��Ϯ�XA�)l`]���QZrG_�&���\/22��n޸�M�*{��[��\F}��Z6 � [��^wu���"�s��ŋ�|��_�b喆�В�v&�wͤ�B���켨������q�t�p��B��r�Y[�+�&S��eľ��"����Μ�} ˜FC�U!�
����j/�UxGHY������vn~ʉC'�s$�rb-+l!���l���b�h]�Ve�-�>��(�/]�|�Ʒ����7(���dt�r{��S��^4�Rnaf�kr	���k���߭��@(�o���Q�e�G�lh(��ߙ�.�9�|��lt����j��6#U�����[����W�d�����Y1y����UYP�=GZEy]B�og~��v��;=�9�&82'I��f�T���@�gKܞR�['����8;�>�����R��Tʱ`=/_�ˢpq?���{��
8;gs���a�Ŝs��� 3�3
��?z��وr�HTn�QÑ��(�w�V�Y�:�l/��0iL��a�Q��L��� �s
43�u����İ=��/�~c'eX�Am�
��(����K��E��r �	`����o?�O6����x��HB�˗��\Dv�"/:.�����<I��ơ�\��҂!������^�.���x+Lb0�&mV�UEWy��!ou0�r�֑��`V(�\}�Ag(Ng]�μ��A�mƓ���~���Ť#M��˯�l�.�;���Ü$.��9�(-(��mx��9�:w:��m����J.]��t�7?B�|�qN�{�i��q��(]�N8�L�s�Qh�릐�K+e��V���_u����SK�P�g��+㋁�?�Ӊ?ʯ�[��&���gi��4�m>n��vgl?�ʭWZe[m��M<J���y��5��^$����ޟ�fkV�B�E����w�Ӄ2����������>hp��Y�zwkB&Qpt0��2߽��pw@e޼\a�>�����sy��C�C�)�X[s�9�r��}��:��ӡ�:(_n[�]�Лf<L�����_<H�u�ͭd��6dړG^���y�=qJ�a��7�2\ui%h��Ӝ�{=�s�[��0�lԧ����h�G��Nӿо��N-f���2@QU�u��`��Ƞ�Pf]Qvۓ[�!lK�;y���}�J�?q�vu�m�F��G��[����6�>]��8y��q�|g���)־�R�s�>�~�}�'�c��Q9w��J�Tƫ4:��c�*e�r��t�r�;c��n�P�J�B�k]���Ч[�lCR�8�nڡ��n��Qp3@uP���/�����*���^骓�0\��,<��C����nA���
��U��6(�e0m��}��_Y�~�ډ���9����~�7yK�e��`R��3�]�����B���9KcШ/�L���>7���x��l��y�ۑ�����/2�(����%���8k����E�����h$"��S�Q����}ʭB�੓K�ڕK���_p[�-� O��a��ަS�#�O,������^_�Df�="N�;��,���
#�Z�5_t�	�|h�`	���.�� H����c���M�u)�{\��˓vr~���Cׯ_k�}��y�s���c0��A�ֽM*f�v��Ϣ��I>�L���lJ��
.X%�F
����s&�x*� �)�W�fQ,'��fY�G��ƀg�=_K����(��ۭ*g��2�!���cFJ��1x#D������ +3��cԣ��ݖ0fn0X�ɨ��o�Ϟ8�?=�y��x��<�ᒈ��^H�>+EQ�����~ko�X���-:	&��!�G��~s�ym�y�� ��A�Pl*�v>~@�ٛʧϽ��N�R��H�y��^7��v;K��ܽ�Pe�s�T�riҶ��[��w�{�a��z��!��lK�R �q��>g������{�k7�0y	����`�J���w��=B%ȴJa�ﱭ�8��2��}�TN(���Z����i�h��dg�<	�Ù3g��ܺ�1���Z���-.��������kͫ�T\�A��ۤ�����͛�\����@vP^�}�@ۼ��mx��(�����a��ep<B��Q����ڗ_|N����gS�ϟ��y��8�����1ao\���;RWW^�d����k��'����/3k$o���_�,-U`n�����v����v���#�y�6r�/�>��G���8��g���{;�7�H[�-yW�ʛ��3q�ﬓ�Ca`�'{���ʂ��|3a�?�*�	��9VzO_xc(�cY���p�t�W�*�t��&��Y;���+2s���
v�+�\�[��?!������ePB�o ��3���2�q�����]��K� 9��[���"�^���U���g/��ȯ7��2������G>RnA�]%���	��o�pb�>����|���]�܃��޺����ᶱ�
�Z���e��+ON�H����"*�o�gy��']o_|�Q�J�<��R���^������Q�s�'���m-�܊}�}��uZ	L]���&n����=sТ�:���i�[2� ��2�1��>�ծ\�L�8�N�aPp�(z�i��jf����l�'�ѣG����i־�/�������9ڽ|�g��A��&���]���*��A�}�I/o��� �8�JVIS�5��g�ϛ��~�-Sʥ|%E.�}J}����s��D��q���Ǖ"��{�WV��Qy\��
v�}���g�����Zb�LW2��R�^1ţN�_JL���ev�/�(m�:Xu
�[����է�w^e�6o_p�y�:KV���Z�9���X�=�Cp�ϟi�����7j�-����G����(���� "D����E����j�[����WT�˲Ό��8n`w����ʚ
��me87l?@sw���d���'=m��
#˧
7�)ipQ!􊱫t<�.{���&>�x6R�����\D��v�Q��Pn̿|�J�Ħ0"ro�K���R9�"�n���p��Wb)�6V�,�H猛���]6wV��Z��������%�2������뙵U��ʎ�������g+����,
��m��D��|f��,Ҋj�Tu.�Ly��	GS.�b���(a��bh�PFz����r�w��#⋗��3�.*4̳.�8�|�_�D2�s9����#'(�6(���r{�N�e�v�=���Aظ�ٽ��N�[����pd�b�a7gl�C�6�/gY�r+���3�*�
s?	\��묋�/�IuL6ȣ�伫��K����=�.G�=�R�`J>�b��i�:�u�C�z@؝,�����D/IF�����ur�iÙg��ʧ�&�^g��ο�=�\?ݽx�
S��{�'7����T��MQ��Vh�2̴�e�����o���)Ĝ�tv� H�z�0⠎�g9ͮ�D�p��=t��\�r�����
�ʫw~���r�bk۷Cؠc�L�!������Rŵ-����cOQ�Tn�ˋ���_|6+,tH�	���n?r�C���O?m�o�N��cK�����Z��� ����Qʑ/F��3i��|���I��Ͽ@�]����ݕ$;�Ͼ������v�xe��7�Y��r0�l�k7��5��,����E���r�A"r����:yC�� ��qȏ��@�jX�2V�u���ш;@�(�E�h�H�n��|�0�,.y����7Vq�rkC��m	p��-�_s���S�����U �V(򍇌�Q�mI�ֵLD=(�␃aȒڳ�lpy�-|W���/.�������%{{��k3W��8��l����v��(���%?䑟i����l�z��qH~銟9���|=���۪�uu�W;�x���+˼��E�:	qû\Q�>��F�t�zx+��dP�{ٮו��=��e���_XeV�}d}<c��^�:���I���1>�n������i����x�k��E=��[���WW>�M�BQ_�+��k�8�
�M�v�ҥug�U��
��?��{��B�/�9���mZz�ջ����j����\tAg�m+�����'�\�}����+�qN�(�W�=�)/f*�%z��@��J��ν�'�m��Z�n8+瘝���6y���t"	jJo��{��1묶#�YYx����4�M*�����܂�A}��l���٫�܎[��P��u�}j}Pd~�&��n���r�Ů&�k���m	����&�� 	��L��P"�Tg�v�2��*��h����?�U��lӚ����^��UpN�v�W����Wg��ܾ�7�4NȦ0ſ�b�X�p��p(���t��e֋���1���Ut��K�׮]i�Q��K:�/?k�}�Y������qs��s:�O�>β���y:C��L%�g�Yĺb�J�4sk��DU��������?�q��?����~ńN���?m�@�����������G?n?���������9����(���:��y} ד}��C 7�{"�=G�ڡ���*a��Jv	��4��7���U{ F�CѫN��dJ��N�W�B˽�gϟ�O���e_����k�s�K�)�3����;�=���a:�����=�^��ݭ(��<�x�(CY@)8�2-
k[�"p���Y���<,�!�|O�������pٵ�Q":���u�vͫږ7k(�vP�9+a}�6�~������jN>�@���v������=m:'G�v���~��w�O����o~����v^tfЯިl�#hswU��H���q2��?�S�V;��oz��t+�
i[��1�3�T�1���ÌTzډ�M�k*N�Ћwg5^elK��t�B���~euՏ��݅�a���q מ��r�����y�����7o!'Χ�qfi�ڡ����ՑKh��"E��_7nޤ�P~V���G��l�G*��ʥ˄��eº?ΎX�ԯ�xu���右
s��iJL:�� c�$��������h�uʎ�%���m:�~�#��j�M;W�U��y�����G�?��Ў�A'������N�8����-��Qgr@����?t����g�I}�	�RƢ����20g�23܈�?	�8�y��t�|����C����z:B�Y�W��m�/A�0� }n�U�r"K(��Rw[Bfn�+*"r��W��5�C��=� �I�
�<~w�{�Ƚ�>����T��$�f����=H�(����s�
��	������[����|���P?�֭&�g�ܟ��O���R��o~�u��/��������Nϻ��%�D)�O�c�������l���2�4|�.E��|��>w��o]��`��$�@[Y�2V�Y���d	�J�}8j��Pw����z�A��<�Iz�o�Ewޕ=�R�2���=�^�:��u��?߾��_<�;���
���~��j&a�����/_��\yɠ�>�-�����
��l�n=�\N}�o7�\nR�u9�6�`��GF���MQ��4p뎲�	�rЉf����N�<}�,q%H? ����n�[]�V6^E�6���Ioh��`������뜅�Q��9�*T��
.g�����°��R8�!��W������d�W٩�ZW��1���ܺů��z]�k��j��>}Y����J�sk�u5���*���_��~*��_���(�]���ۘ0��CA�b�:�j��qF�{<�0�ui㫯��֯H��LYf��8�M�]� �ܽ�}��F;���r}ZU�ͨ`�4����ps�~��F#wo��s����+,`��:��l�B�׃\�}q�<͌-��DԴ����ȓ���e��B\a�lhU.;�jF:T���r�3���|���(x5k+���+��	���W�U��U������<�r�(m�!�3t^m�|���Y�v�O��Q?Ŵ�C`)��O��)a�G !�+5���y�'ޥ��D�knq��fj� ,���.�x(g1�;!��K];�:����Η�B��a�%��湸x�����[g�=�(
蹗��Ro+p&�Ω�t��Kq�-�af#��
,x�;�U��P�7Q�v�Z����jm�/��9jV�u���\�V)q��CbPasP�v���Z����w�W_}�~��_D�/��k�楚��=�\{���{���u6�6K�5X0�,�Y�)Q8��@:�V����9a,���O���kݻ1�0�1↿�^>T�k�,u΅�8��vW|�R�^�WY�q��:w�����}���]�L�D��:m��I:C%�܂��<S)�cV��8��~�v{�]�~��'�����2@Ry��(ǟ�2�*q\!�mϟ��=A9TQ��T��3����T�E�Wn�R�P~Xg�L��b��Ƿ�.�J�[N�S᳍l��#�5|B:�Q~]�q/�c����
�%sgy\�<QJ`,;�'�Px28��$�v��j=���;;c=��l�i7%��+�3��]EF��$l�Y��f�t/
�B3��I3�]<֓��f^��AG鶄�ܖr��ʭ[�\�[~���d����ʚK�(������K���}U(\�u�Q��Zs斾�v��}Tn��@ʶZ3]�ɶM' �ԝ�R6g�>p��
�%凝�y�
���(�~�>�w��o����z��O��W.����-�ʎ�?�_����
�@>�����M�����J�&?}�x���4ׄTx�g2��$�ď
�K�G�Z�R[z�uS��쭻�i %��$�����7W��z�^yW���~���ӹ���1�*g0�Q�ABp&ЭH^ͩ"��)�^���vݯ��h}���L���u�n����y�{�>�4����P@�,S��~�O>���4����T����~h��sY�G��v��#V6<Q�ԕ�ϟ��F���=>?�q@�t�e�����h�[]��$[����[/(����N%WY �L���Uߠ�n�W+�Qf�K�b��'��urOQn���up��X�cc��i�](�m�S�w&�������K���������I;��l-�d�	�$n ��(��d%�r�'�j����c���̋��Z
`g<�8�Ќ�N%���̲��گ���}s�������FPP�,�C9y05/%� `d��7���(��&�F,#!���#(�m���l���GƖ�FM�}�zr��=]�R��8uu�V��S\3c[Za[w/�4��4���)��{�n�C;{v�?��p��{n�{��p��B���=���Q��58�k@�itx�/�J���ޝZW�����GS�W��$�1t���uӉ�q�g�1�.R���ѫ~
�K��
��k?��*����v����=9
��;˺G�Fe'K6����c?9H�oT)Aʤ 6;%;��eⳳ�����]g�i�uY]��H\�٫�L�Iᓙ��|.u��z5ٚ�o�Tj�P��C�:FxO���W�d�+�K�ݠPc�
�[^ٳ��Lܥ�3����A޽w�}��7���;_1�V�;��ݾ�A�[{l��Q�=�[gn_�-�v�����u�}��˪J[��=�+b�_�c�.�� @�u��?�'�k�?��f����;�}�t~�F��g~�I�Ik��Uˑ���)rƛ0�#w�<hw��7P<�Y�0�Ͻ�����PHeM���D�XR���w�..�m}���G�L�Ϭ��/�lW��� 87��Yc;�;w�E.��s�����Τ�O�svdV|��id���^t��Y⣤ߐ1]���^B���P����Si�Nndv�7�C|�Z;od%e���_ t���U{��ۣt�(it�ߢ��GEH�z8������jw�?ow�B��&�W�IW�(i��_ꋚ��X�C�L�|��{)��~S/���U��e��A�&]K�ڱ�����m�æx5���j~mi���5P*���ߤܢd�"��`��h���Q�UE�~Q���#g��)�����U�(���S%W��뜄�lIWRp�ᱱ���+=t�`��Aʍ\UH]{U��~p��*��6��y� V�cc�w�}���QL�D�3o��o{������"Ù�v�Rf'�c�g��J�e��'��s۪}�3���a6kE�����T��ՎB�R�����*�t�٧2��x��b�3��T��s8"tSf83}(�q�Xmu�+A?���Ѯ<,�d���^%j_l�k�׳��?�'�?�V\@\����UT�ph@���n�z��2�I�Ͷ���ST	.\�n�f��~iԳ��ʒ��_�/8��~�Z��	�~���yn�q���~��Aˍ=�[e�"Q
�K�:��p����n;S���uU��`��q��{��)_r�09PϠ|�:����:���n?x�\Q����18x+BnR���g�.�����#����V,2���%��`}�'���֧z�[SQn�f)�9э��ό�J��EbIBr�mb*�V�3�Z2�
��G�*~���jVP]��(�\%�pvJ������^>_k�tN�۹T���T���O/0�=|]]��~�8;wB2��)�Ii\~�֓�΀����6�@�_�,���q�N�����9���=V>��AY5��Zh�Еn4lg��u�3gP��eVƽ5"��V�d�\�ݝ�A te�x A�JH��T�^��y^�ٝΕ���+���X���bAX#4��eh�(!�,� �O*z��b��s����l����[7��=��c _�WG�vj�t�j�/��@�?�@���+���ѧB=B�N�!�K9.��Ԗr�Qn��ޑ�S�֏3�q*`r���z(�]�s�c��+�r��!o.Pu����A p�eıϩ�����F;�GLr����k)uX�����ҙI_;q9�ox;���f�+b��˗2��v�;8�ޝ���=+��KM�^%��/�5p����.	�e��,i{�}ʏgm\��y����d5�
�t�sٵjc�Ξ�eEW���_=���eO�|��U�l;�}�v�� V����ub�g�͙�̂>KR
UIe��~gI�^��ˀ�18�YY�C)p��2����ݷw��<�� �8Ub:C�~x�R?��оv�f�u�4�衕7�{f'%>�����폚דIc������$/�[3ع�r�)a�76���(�u-tP�����Cv���!�% � um�A��J}a������lnEP��J�#?����8�L�%�b��;w���N�����*�U9�)��t����9A~�G}�<w��Fi�Գ}:�0�%��t����!��������K�]�;��~O�X�m�2�D<:e�78��L��ӯw���Q�F셒��i�g���p�쒎7��1�c���a\b���Uv�\}��T�W��W����]u����s>e	�7Sn_�oPޟ>|O �>��V���M��:�W��LE�/J櫢�Pbi_먾�����>!�¢2��o���C�9ȟ���3�)�������R�g�y�*v����.T�SJ�+1�qW=�O���{�B��\�a]�]�S䫢����C�$q�n$8~�E�߮mj��8#�������(���X��|'u]�K_������(���ʃ�n���Z� ��[qx�5���~� ���/^3��X{\-smW@y6yR>�n[��҇6Qb��`�ȉ�u�V�����P��되�\���vx�|s��)�_`U�vB4���[�Z�v�%N⹽��zA�i�c�� <��<;!�������SpD��k�q��U��IG ̈́��aJb<���l�v����^���{�����(���\O��o�ʭ�aq���<�N�옳�
nJ1�ڠ�p�3���9u]3~�wY��Q|��eK������OaO�?Cy}��]~.}��g�U�V)=kw�<��W����Z����Q;�E�۠�<�bc�*;ZX���Uy~F]�p�̚��{�'P<<�+����J�5:&���uߨ�Wu��'c�W�bVpJ�J��3rd�@�X��N�
/�Fډ�OO �{�Z����Q��)�EO��㛔	Ƈ�_�����Y�ѷ)�+ ����^��}i��r�u��P�<�a[�⁐����z�}�8�����^��-�[@T3�5N3S��Lg�<���B�CPj����=�y��dJ�A�h��-ה\8�;��t0n?1�K�.Ԛ�w�߃W�>u�D;w�L���FYr;K�fB��=ׇ���-��[�疶v^K	J֥_�I�;��N]�g�P������O�,���bb�瘽��o�����/�],}N�*�{�{�,�6B��;�܅��MdY��k�T��z�R�MZ9���׽k��� ��%4:��UD��T�t��K�N���9�D'�~g�7>i�|s'��_�;�\�~�-�<ְcpf�>��$����W�������@��̼;󶼶�`��v�z�Pea��\���HO���g�ܞ?e�et9+b�=%!2p�绻�3�����s�Te+2����K��	NDx����e@Vֆ|�����U㣞{�W��V��
���<�$�d���ݗ��nfi�����������*�K���=�_x��\[:��"�Z��~��g�2�E���yR���쬠�>��û�7m�g��þ��A�W}��D&3z��	��|.�֡"g�vIG�������+/Q$U�ꊻ��_�Y6eйv�����g����۷�-��ڻ�"��!O?G	��G��߈�{���v�*�-���|������Ń�>�R�F��3î���O�ћ��?)c�$z~z�����7�d�$�QVͭ)(\�(<�/w���>�����󮀳����Y��l�ֿ�o}[%�>��ag���������܆G���r�9������@�A^�����r�&��B�kEB��AP�]�xm/�(�*�N�8���QUP�Nl���"["hӱ�W�h�w��{&��������Tj�:β*��se�����TC��_�;��f��;�=����Џ���'Jr�v+�3	��8�� @[���+�<�-�BJ��5ѳ(�W�����w�?B�x�~9C��(��岯G�#�0^��>7?�,�煼.ë�k��J�2'�\&|���qr�2�������!�|
�����+䪈��N��^Ľ@�r�Ϲ�QT���x��_R�8"�<p&#t�a�o�*/�=I=+�iy�����������9G]�c�'4���*g�TX�jȥ.g1Ou���R�j��
=�����)��23G�2|1r�Q�3�BќQw��SJ�^3
A��(���S���V�F�FV����1�+C"�*����%�����#���2/{�N/�,���0
�3�uѽ�m������A~:ґ�붱�r���m	.%�.���Ah/�?��Oڿ����������v�|U�W�Fp;˷�4^�B�+�C����.]�	K⁽�iEy�� �87��^ܚP2;3��T�SC��p.1��\<�2��������.�@[:,gc�yu�!~`��3�v�P�[[�-A�V�zm�����_��h��nep9z+���m����|`9Ӂ��h�#U����UTjDƶ<�x�>AR�3=��G{�!�/�x��I�:�t���x�;懬'h�,8m���O�U�Sձ�T�P�c��(Q�����(��*���6-Wl�8�-����r �ܻ��|�6g��2r��;�g��O����3(��[��+�nܺ��s�N�E��?�U����~��_�#��O��}��g9q����������=o'N-5���'��O�u
i�%���?�y��/~վ��+��b�+������v��Ep_��yӾ��^�������o�	~^�������!�si�fƐ��̢���z�V8�*�PjPd\�.o�x@8@~��j_>K��Y.i�\�6�f�1�p*P�����Ӷ�v�ɘY7�?ރ��
yG�n���������+"����h�ƿ�?��g��)۸�������lc~z��M�I�2�^Рo���U;�Lڦ�c���+�N��ᇺ�݃���9i�o�o^{p�np6�$�c�msHr�L��<�S��	�D�U����?����O�2��Q���^�i�����������o�:�ȫ:��?�ۗ?��n�:�N�<��5��(����.�d'~Q��*����F�ꛧ�����YJw�Oz���=�F�I�"!0���H=Ņ,�+w�q�F0h̀���C�;[�����M'0rG84v��}��7���י:�m_�-'��(`*�*���+q;���U�C�q�/oK�M�|��f���2�n)l�{����@��j����f���qH���ØV�A�Ӱm�*���mU:W���4��	vB^�1ƏݸU��eW�Or#͚��8�Q��#�/��`��uP��f��/j���,����+����]i(�J,�$���z��W���~����Rn���I�G(E^�1�ۚJ��M�
x�F�QQ�� "3lH�N�a���^aE�C�R�˥R�z!윦�n���bw�U
�@]�/x����4D�H$��R�IGf� tta��[��eK5����;j����*l*=�S	K���iFɝhTy�ב���\��r���C�P�0��rK�t�v6Q�M��,������޼F�5�Aċz��]��?�Ū0�1K�>��3�2�Q��[�c�J�D� ��t=i\Qt)�ydf�t��-��Г�GUvk_���ԯb�㲘K�ΐ����N�db#;J��f��Q��n{���v;w�h�ї�ڿ���J�C�۫�O��Ah娖zt�����bE�SeQ���i�p�2��~��o�/�}�
��/�x7�@i���,�u��e�yM�6e\l�>���:
���ک~
U%��eVy`#2�C��@��W��P;��r�6�����?k�r��7��j(L�oe�� �[8��RN��d.Ey�K�O��X��_���K�%lO$6PY��&��t�8�������YU*�f<J��O�ɡ܆'M#�
��{�A���ɠ��H<$j�^�n:�/r�:Ad�G^�>���ݒ*��uk�ʭ˾Ϟ2�A�Y�Y���?��vV�T�W���s�ݿ/r��G7���"����=y�����U�D����t<��薜������G� ?����Y��1����/0=E��=��HS��B��rו2�W:��í5�V�m�-3l��g�x�#�}m�f��!N�@�?�V�[yo�1Y~p7��1������؟�t����#I�h2�}�����>�~������]���>%_Rbp�$�3���L��a���/�3q�`W���4��̽�_�}��������wW�����ߖ�d0it!��'�2A����1��MO�w�bx�O��9�MeۗZ֏�|v;�a��g?�_o7ʡk�9\Yy�|������ۯ~�u[Y_k�ϝm��?i�~�I�׺��,�Վ�IA��*�)�f<r����A���Q��o?�3�����C��r�r�M+'�m+��j���3�1};�a�|��(�K>:�Z:W���|��mܙ]W����!&W�=���X�( � ��Ӝ����Y���A��5�����[�0�bw�����V:�W��7��5X��C&�|��ľ������=-׌�w�������K>��<uP�,��4���s��!^�MYIHe_&�J�p�����k����Mʩ�A��|�O�� #�2�rk����V1,��!�� @����3�����r��wPnf�֥1?w���ĬD��I�Y(G'V��b�}G�K�����"Ŗ��+<��I�`g�d�Ƽ��i��b�jƈb B�B����c�agH�
�����y��ť�Au��ď���sj5 �Kh�t搉�]�Y��O��/i8k$S�@�8@C�j���[32� ��iJl)ٝ�Oj�S)F��(Ґ|�)�>�q$m����#lR��P묖�Q4i|��h��������ˎ�${�9��tgݜA�C�ϸ��}��_u��YUO��6g�lޅ|���DgI�zw���%�[����>�����/�?P��z.�\tkB�&�b�O��F����gTi�'�S�l�����ߠ<~�~��_7oy�ƎKw�-4K#$�D�~�xt8Q�?�>��F�яo����4�K(����}��@~����+∋l�%�����3�?o���۷�>d��Վ.��z �2�����=tɣT��>���������{��g|�;o����0�'+�K���F��[
�V�F�)�V��>��BgR+.������{�ڃ?���&a<��'k��M+�:���r��m��/{"�;A��|���m�{=s��e:1�۫ݎgI���MloyG�_|�^�x�
?���^�׭���C�����'D�x�˙S�2�%�s�V���s���������"����v�m�n�n��嵬���Pa�=�Zso�|+�̬+���Ç�)K�l���̄�_���<��U��k�3a+��q����6����ߙ!?I��׈1�������$e����jwۏ<�k��d����i�����j)�g���c�6����)"�49i ���QF�-Y mUp뀍[䜹�G��헿��}�����_k$l:{h�b���.)��W�kO!�<�����?����ʥsԏ���F�5��Z2�D��ށ}�##N*�W�W�m��ߴ_���'���~��ڋW��"|�ٗ_��7o�g}+�ۃ���..� ݾp}U���m�a�](z��W_}�r���J�����5U�����������.`Y�M�O֒�ucc �����	�J(��-(G���'��9Q�7a�O�E	��u0��XE����@����)/���˶h���:��s�xȝ�[~˶�D��ҋh���68g���Y��t���C��v�+�E�J�x��J&<;ɗn������Ǒ�a�ʞ�nZ�����n���E9mc�}VA=�^�̑~W�l#ʖ�����ٲL��CBO��?�r�:n\��U`��O�)���4��Hf�	���9*M<�IX�B�*
��V��
RD��o	+��E��'*e�Fn$�P��L�I��D෧'�1�ܐ]3�j$�}?0u6R�PYN��q��`t�P\+���%�RzS� xFANҤ�j8��k{A��ŭ���=ʐ��I�^R&g���қ���� z�D��ʗ�$�� i7�WB������xZ�M:�T�o�����k�����2��L��+�����x����V�ۚ��םep�e����䖑Z�7�h��*흼j��t����U-��V��R��Ȁ(�q�ϼ�>��ı~ܣ���=��wϑuh}�V�)��#�;�B�q a�~`o��7�F�3�����A�
�S�Bw���l�/��"����~���?Yɾk��{��U��j����%�����T=��������_	^�1�����`f/Q�Ҍ���O�#��OBR��݄�yO�d��l'�.�tm���fYvc{q ���(�<�Qx7�`�G��ʰ�Yj۪*~y@��3�2�;�sO���=��!�5���0�2�l�X��ms�R�셳�S��C��s���p��mR٧�_p7?�Qf����M;���G��,��L��,��sÇ�׵B�@2�+���`��tF��/��GmY�-k�M���)��H�:4�Y/�T}��x�ǭ[�4���$C�3�POK9;�^��a�+�[��Ԍ�w�޾�q�zFo���q��T��&d��r���mh�n=[�M޺Q7��qgm��yt`����g`�#`�1��u���cy�}���Q����0X�ڮ\;���O'��^w��A�1� z­_'��.x�[����2���VVߴ��=�x�y�M|��յ����bw���(�+��m���E�����~߾����|��{�_�ȣl̹���]W�.��)��� mպ��Ǥ��P�T�i�򟲳d��k��2Ez�� ��������:�i8�S���g�L_a�u&ɕ��h�=�i�L2_�]Zˋ��:��_ր����t�AN�igV�0�˻�	F�ҩ|)t	yg���a�a�ӻ���Vm�4�8��:������F�����)�Ƴu8L=M�Z��2ֳϽ}��䵃4����%i����%�P��~�A�\s�"a,	���-eӜ���I�
�/ʌ��5èC�%z�mF<#���K�h��z^��D��Z����%yҤ�����O�d-?�P����O�qH�Rl,C�4�`��lƑ)Ea�K{�7�L��均���S%ѝ<��m=[.Ört��@"����+K}�Z 1BR�'�11i�(��KqM�{e���#�
��`�x�����4��P�ЫȻG)'�#��叺R���f�����Yf߽���s�*���U<���?��
a�-���w7��÷Lg��r`�Uom𓚹��|�Wg�{�%�^�O�ξ��mk^�C'��NnG����kXr�;8�r�J��N[Y�t1��.�����ث;�_Fyy��A�����:�'�O/�P�!������[���e�V�[���-囹�lA�N��M�Ra��x=����2��ϗ�)����|��)H�����|���L-鑏u�|�������ދ7��]�8��ZrsV�Ctp�,ŏ<��2��c��zV�#$H�D����RH��r'�y���nB�R�s����>N�Wy!�QD����CH3K��O��"�x��V\!�ڲ��<�� I�
��bI���e�1+T�0�Dd�F��Bc�y�����LO�~1�ǲ�"ʹ��_�<��w�)�j��'�ݓ�MW)���I@<�T�����C9��ɉ�M>�3Pu��CL���So}y����.�z;���PnS�e���2u��[1�]8��_<Վ-)K�N�gy�q�rfV8��|���
�;X�s�N,����'���7�g/3s�G���!C���W7Q���-��v��G�H�{�[6�f�R����yx�����X'���*����@��;��ˍ�C�Y��6�-��W�g��!�N؁�m��T�]m��Ld�^mu���jC5�RyOx*���L��O���`z�k���|�r����C�<�@�2c��Y�c�Y\���I��Jw�<{���i��=2TY�3nU~�	�k3w���
V �b�[�~1�e�k��>#�����m��f��o�/�����[?K�BH+na���j��:>KL2����5�ף#�Ô�?��4�t�0 a�t4��i�4�,�m�G|���h�v(^B\3<X0=#T`L%@��4�-��Ж{^I/F�ٚ0dp3��e��J9�������-�$��`�ȟ~�cC*b�.��LL?�� !�O/Ao�vj��ǰ�;|�.��R�卩1����s�=������"
l��c y�Y3p' NU�E6�!�*�Fc���-�q������t�]�p:w/:�rƻM�-P�	o鈩AǏ���w�Zn�%��J��B_��%���avZҠ�?Q�R�q�exC't��=*�%x/��3��,���-�{�Tp2�SR��i��zhD�.om{!�_|��K��˧�7=xH��tK�4)� ��2=Jׄy��n0U5�ڀ�/�J�3Q�"��Ѯ��e��������Ί�,�Q��Ey�t�Y��M?6�M�:_���_��rgPd�e����y���#�XcP>��|�g�҉�6�s�,���o���|�'X���p�n�s�:��hɟ�	�è��яIH��P^3sJo�z����m&A?ۈ�L�����I�Y��,˻mǭL�_��D�XV�$��
��|�0�N��gka���t|���� �[9'@�MIr������ �ݴR�g_&i����(��/h��]ǭ�������ƍ�m�䉣9d�a�l�W���L������� �L: �`)G<e��	��������V��P�FN˓���(���B��?���xۊ_��2�z�I�|̒{�z7�y�v*�`9�~�MS�;��<x��=�%x73�nY�J*��P�W�^\�p�]훶�r9�sܺQ��Ƀ�4���s���)O
$i��o�Ů0Ԉ���� �6�{�a�AM�h���|�_��Z �R2V)�=;�]:y��ʠ��Q>�H���(��uކ7��M���'ʙ����1��]���N8&!S���бS��d4q����廿⠼��"���S��=�5>�Q�r/G��M<��&����o*��l\b�^I���d&UE��⻻�Iy=ϳ�Ν9����o���7����7�3�ZRj�綾��pL�ɦ*T&���3�U�0>bF=�'�7LwK��=\�5�G�X����FN2��F�9J�M�zx�� ��0��L�f�ƉS�ɿ��5�z������y�ɐ��x�����kX�y��%���/���̎Ω�b�j�=q;�8*g�����"H�\;av:k���-�c�8�=/)W�|�@A�]d��rt!QB���n&`8y�� �!���m�n}���Ndyn1{��pܓ����/����N���� a�>hgW�L�$8ۖ�_�Y���9W�<�>�8�F����K�?i�2U
��v��MxPȯ���
�;
�&r���8�u��k��qÎxɯ��2l�xQ�6��$���}�1=�4��m�x��S�k|��Q�0҈�W}J�z�r��p��zGk􊗈Ik�1�e�w�{m�)�N�+�Kɘ�5 S!���	���45�̷��0����_���i�M�j�$�(5�5��`k������G]�s��0�gw����n��NyM��bڔ���Rn���zX}��n(��iy̃���<aUl�)h�G��D&��WcK�jC�h�K�I���������ԙ��Aٶ��P&�����귘D�tc��?���%S�M�rV�/�,m.-z�K��� �m�	�З<�U�z�t���C�P�R�2�K9(�5J���R���'O�<�F@d x�l��h�9x?��s�څKgs �Yf�+�g�[�?m��Aڔ+�Π�<�+���#�lUW9������:�b���}��C�%���y�
��v��b��`]�����40�+�������M#v��H�Wԭ�E��~d@xzz�T��U�l;tӐ2w��]�Đ�Y�:N#��\�x������pYE���������t����S~#)����khJy��W���z�~�g��,�Y�� �C`�"t�ӌ�縏��ń��m��5�����'�^ŵǿ��e�I路�O�:���n�h����΁2�[�'��Ch�G���*��a���j��r[�d����%�T��3�5�m��y���������8I0[�H)��W��J�t;A�44�3)>��af��0o*�x�*q�}��xW�������V�u��b����Y�pgܮ�!z�rB"!�f
nf��������T�g�t���T�ђ�
'O�Ю��~	��(�
q����O�*M�/�>+�l�t��5KOpfy��xL���bP�C	g��go2���y��-�Y0�ޒ�C�d���fF�2I��'���!�����#��t(C�7��K��8��4�[�X��$��0��$����B)����j�n�<��x%��l���?e,s�ې��^P����F������J����7�q�(ʭt��Ho���Un�1��v��Dp��BL���O����ڍe~�9��ܚtԴgn-k�ܢتܢ�FaQ��A�ց̼r�L�~3s�R������ܪA����L�yJ?�j�34� ��{v��&�o�]��j�,Om����(p�<J�b�'s0��5i�>~#8&sd�F�k��"�օ�lȃ�f��~�_������	�޶#����i�I=����xd�_���Va�����#Ȑڟ)�XUxg��	G��\��RK�ĠN및[��ʦ�l����ZE ��Lt��yj�� �;Q(��N;�ww�����r�y�B�ӑ��wU�{��,@
&C^��q�,���H�J�R������;a,ۻ�mOkz׌g�a�aHÿ�5��mA^�M����G��l'��*�����޴���I�5���>ǘ.�S�Vq�]�f
^�{��1�e$�(�g��p�}����q)z���n�wl~�}*�^��`@����4��a�k��}Jc����\����Яh���n�pr��F�}������*����������c��"K'��C��Z�.ʐ6Uf��Զ�Un殱���S*��
����_���ܟRI��y�ϧt��X �:�zU\S�ʚ��91	W(�S��(idSOF�)a���G<��y5�'\7��R�����g�q��T�M�{Y5)1��A��+-֡e�$�LM�PpQ8�PA_Ïd�Ka|�BTOiR�H��hV��-��rkZ�5�4�?���O�F:>k��
��u����Q�T.05�b��E0H;������̘��݃WBV|�g���km���4�ԓz�&yVy)e���PӁ,G�[8J�Ѕ|��ټ�#�6�3Q�_�����*y*8u�����7�?�RALj���F�M��FH���#���u'�3��N�╼ ���ߘ�����R�d��ڙ�d[��E���Dh 6f����az��&��'�p�\*�����*�(�;�[�=������[g�I.�r���-A���Tn��ʭy��2�ڹ�gmھ��Sg4P�3�[m�d�7�y��i�.o���j������6�s��M�L�h��`y���F^2�>��z�}�{��4��]�Oٵ�v��/�}"䇮�Q�i7�=���À��M;��b��$�4KhPA��G��Tn�d`�uM�+��]��^�{�Q<�V���o|�zEԇ�|8��#�Or�(���p������,���{�֬��_{����z��=A��\Jֈ'�&~3��>o���R�f�ڕ9}b,�ۚ�2^��M�Cp�JR���K���X=��̧����<��H�|�g�b���qI����H'��@j*���4)���CeQ�TiͿ�&��6�Ǩ��2gt ���嶃&vw�1X6�M$�e��(�M��ЛRn?�����Ɂ2?����<$AOK��#�����R3��m�!L�@�\��H�\��R
L@A1g��2�c�0�@�� ҠtӶ����-�sy��N�҅r��ki�=�Gݽ���}��L��{����)�<�'?sP��A9�W��0gfoUF��VF&��`�w�r�!�#����wR��۸|�Ğ�\ϳz�x`���}�G�{�x���ħW&y������:�U�m>���Ir���ލx,ϵ',U�P����(o	'o���	�|�ý]@}��/֡���[��!��l�Ƴ��yY�������Q��7?�s7����{?ǣ�Ln3S�ӹ�:�Y��Y�(0�&+�%�����x:�m��RH�4�a�3�<���t5���j�����?p����3��s�)�ࣃu5��La|}z�eЧҋ�E��⚧~nS��@Y����2?��<=x)�?� b.	T)ŉzJ>��ݑ���m�y��nE�z.���;ջV��c�$3{�a������ELb%k�]4����w�ɇzR�U!TA��[�3u�K�7K�� ��m9i\��:*yg�x@�c�j@'?_�Om�(��xȯ(:����;(�[os��ζ�Tܖ��f�l��L�I&����j�v��C�58�>S��b�J�~�}��G�@�,f�t{�cX������ s0=�}#}�%��e��7�Q7���f�
V��Hk�y�zJ����p#~O����7��s�ן��9�uWy��mX�u��̻4�+���^y�<������E�L)v��g墼3�O����i_�ݡ�ƻ��.�/���5HA��v�sgO+{G#!FG�`F��غ��O�F���ڪ3R ��"�'8�/R����Cq�Ӏ�5!���������m�0Py�A5%�����t�r��]V����=-Q;�̹�V3����\����K(��un�{�(�,o��h��U���
�k�e0g�Ay��3�nU�^j.� ���ǯ�}0GG2������aK��Ӏ� ʒ���*�	PTPX����j����(�(����uG��������[:��8�y�
/���������y"��K��L;�v�뺔 ����v53���m�;�3�B&��v��1��af���Cf_z	��x�t��*�R&w����H�=��Ow�P��<�Ug)����#�{�P;���3�f���.c�b�yd�l{�7�'�6�V��]��{�˲��tN>������v��\�ӓ*$�{�������c�en>��;09���C��{�c�Si��&q�5� ��"�j|�h���u��YOe�¯+�����:f\�O/C��g`�X�O���ӎ�TNߠ�<��E�#L)�~}���𬫱�P��*�P��u%9����e�M%���K�n,�$�F���o��5��$�e��}5fZ��od�K�f����4��~����}�ѯ�G��F�P󃐏�(�[�+ΐ�w�<hx�;/N��W�獮�Vř�)y�>	�n�Q�`�\Z�DW�G�O� �$_�ظ��;�8~���E�U�C�o�;?�S�O��h~VN�5Rfn͠�DL�Jh�Ԇ���,���Ry��l�Rx�m��<��e�,��.��s~�Ւ�G � ���aG@�N5�z�]���*n����z�&w~��?��Q3�b���Yw�Y3޻��1���<��}f���ؖ���Ŧw-�S��,����c�o���20[
�;�*R=��&&���~@�;�)��<�֡�ǯ�����ݬ����*6�نA����<��Mf�"����D�D��J�5�^3kv>�e#�j��W_hK(��&/x����& ����a];�L]aS*����<D�e��0���q��Nbǭ��Gkv��a;h�M��<���g7��OfnӀG�R.���1���`X?���)�0Q@�l��R_?.�����pqv=O� .�4 ��kf�2Y����)�~}0FL�)�
�rW��t?�<耪��$?i��A��#t0jOCo�=���U��+^�����l�8��'�I�{�}@w��Ǥ���t�g�o��x�`�$;܌�a"#?W�g3�ҩ��A�I-lz>�h�~�9ኌ�*ծ����Y�q��Z!�z/�3\F��%c����1��ǎ�@ƨ��/�+D�q�������"c��wp����cO~���<y������pw������ׁC��jC��o��<�[fV���eL����#בּ=�5vx��7L坧=�1�I��#힆���Y߼��T��?��MnZ��������K���̬�e|��p��F��4jv����>�7�5�����Q��ǜ���'�p�M�ř[�o>w�T(i�ʯg�7��7i��Trq	*����u2���ň�4��d���������޴�GZ�c�5���/	y��+q�dE��ߎo�)�,����PQ�(h	c��n��C����a�̞0���O���1C�j��@�� �Yt[�<{��P�P	�ʝ<`#����KS�c�̺h�<zڕ�~ ���>gz&O����`T���Jp�g�a�����8]q�A�/%S�W)�N�e��V&��t�����gv%fx ?�s�ݭ�YhI�Qs� ,@ӿ���3�{���/���$O��&�$���p~�;fd�6��*=z�3Ǚ1�ЦJ�=�D'�9r�f��~� ��̬j�h��՚U-����}��{��<)����{�W�8]!N[
%��=4��*�x�7���%���a��V.}S����R�t������T���{���=�������f��~3y�P/��~f�_�䱗��C�Y?����P<J6�Sm7����k�˖j�R��s��Ϳ�*q� ��tЭ�MR�"32K:�%9d���AU.w\��=��'m�m����vʶ_�]�\���}�����V�:���[�QJ�t&|���u f�(C�����߅n��4ELk�͹�������k��5�=_��u�Q�c��!��Aff�=��޸�}��,�����n嘷�Z0d��򅲤^կ���=P�v�sVfM�˟��GF�p��{A�c��p�R3�C�o�/~�%�O�>o�kj3�x�1GrfLr@ޭ�B<�R�m(�4�>��d4t��3p��v?�O�y�Jly�J�v��v^��U,h�~K}4���9�\
�Q��Z���)~Y%�{<�Aj���8yi��`���遦ps��3�7L/�~O3�V��MB�q�h�k�s��8�>=�6�߈��!�3�ǘN��ZŤ��i�����G�Oi�^��/�z��wW�����<�Ʀ�o�$�D𖝿�p}�C�$(�-U��T����A��O�t�؉k�J7�D��y�xa�� ��I:��Q��}o���@�L;�������ߜ[2���T���d���7U��F�1���t�������u?�e"q0�*�*��Q? ʯ�vɳ�G���M+
oWv}������E�T,)�ex��mx�J��R���U�ʟ��q����A�<Q�)w�#8�u�tU �jJ��4SF�8L����N� i��GL�O��ݵfa�p���{h=G�^/x��>3���j�sާ���KhcG�����6���TH@�&?ʝ>��Nک�QwҸ?KO���fփ�O�d�K �r+R��u]�ry����_X�< �+cT>��KP	���2U�%��Ė��=�B=)��y��Rv��nlQ7ɛCn$^�g1�Lu�K١�������%pu"meVg$4��t���Q^L{�v�W����6]���)�R����̥w���x�{y']p�Jv�:�@���
)[��՟;�4=�����I`�&���#���.<��P	ĭ�"���v[H���ǖ�E���[�=m��R�]az�z��4��myH٩��f���Ņv��I�ۿ鶄���ً�܊�#<�[2��iLڡ�`!�@�}��
�lmm�-e�J�R{Te���x�o�/�E�69V��)�£�y���ϸ/�)�!t'�ADan��`�A8Ml��!�?�����q����0����̻.e�/jF��q���y� �}o�E�0�;�_�;;���ξ^xG0��V�<'ݎ��y�`��$Z��>�Nz��p�b��N}�����v	w� g� ��+�.�J;�fgw+q^#أ�8�KiHS�
�!�b��(�Vf[i��:�Ao���+�:vՁ���`�����*���a���?E�g���Y���_&�j���$�0xg/T����0�^+�;3�[�u�R��̩�I	��ƕNE)�!P�<}���QK��.��g��A7������'�rӬ�X�)vV0d���;񢐊kE�jٖ�F���S&J*NQ����3�kÒDڟIV��DZG�%�	�n}��|A;�ĒF�IZ=7�{~S�D����]�A�S�v��X��|	��9S�gy�L�)ML]�7ä��]��,(Ţ����0�q��ئ�m�ٞ�+%[��(�yH]N�$΀������öX�E�G�����ئ�������.ʝ.s���Pp'P��>�s�!-���������O'<~�e��E��=�@�`���	*^A��P,⃉
�t��8�Zt.�������ƻ�- ��1]�NS���?w����x}��wM�)3�W��^\'7�{�2oH�0Svf�4z��^�yV�3����]�V)����2�Z6�i���}��)�y`؟Z3;q�w�_ݖ0Sn_��[��zR��f^��!�@�����Z(�[?I��V�v��� J�J�(�~"m��� r|�X�]6����������/6n*���:���O��_�B��N��ц�?��C��h�X2X't�kǻxjތ�)�0=ĭ�s��u��Q��'>��I<"�I���uW��T9cz�s��K��׉��)i�n��d�[�1�aƥ/���6�d�6���I/�1��q�S���J*��o�A?f��Y
o���kf;������vx�bd�w:���hE\������,-M��%�|��|߼�6[�iG^�#�����g�C)�Ca�Ď���u����s��p覓�� Ր���_�ƤS�̻�����c���af�V}ό�S;�՚���hP�y��V����v�����>�}`Z�yr։�oP.;�\�eG?)�ԉJi�0T��|�c���{�i�ٶ ��[c)9F��s�\RPy�$���-[�؃�S;����g���a�E��͵����afa��`&~�♏��3��a��}���wLxez��m��V�u�m�)m�Y���>�ց �Qo�q�l���}Rm�d��3UA����8�;̴�[07�+*L�K�f�!7��H�ه����k��2�+Ų�Z�O��
*����"���|�*[xNG��V��ɮ��?��w�1F�R`�A�xj����.Mff$1�t���63����9�F\�rW�3��A'Sq*���e<ۯ�������_�q�Ëy�w�f�y������-����x�]%���.�r�Z�ﱏ
��;�IGQ�w2�?����C��Ъ�n��<jG&���������B;�r���[���e���=P���Xj�	T���@أP|��Qj��.d-��1gg�c(�*��О�/Tn󼸄"�B[P�C�] ����!+hL.9z���Ȼ��9�	e&�ʥ=���������M��ާt�~���c�xfQ�����S��:�����;I�`<l��0�4hTI�7�
Wϳ'�'�8t����0�/�b�=�O}h��:���GX�)��6�΋���b����L[`��R[]�-F?��u�F	�
.��WG�ݣ��.�_/�O��������E�|�0�7��- ���}�����2"���[t*tHtV�k?H����sM�f��N���<�C7	�S7L���[�-Õ,覻�l���5ʒ��_	I����?�ݣCյ�<gJA)�n�cqMl�33�����1��n�Ҫ�Ԍ��i)�v�>g�UE�ʽ��KG�`;{Ӌr[�|��Dɰc���̭郛��jF%��)�=��
sU��4S�{������s������c���}��*|��7�7��o*���2�34�x��H�S�����QcP�����γuY<�����75m]۶�vo)_
��E1`@��÷'�����3��Û�,eu�Ø��4��	g�C�����Q�MG~2:tO;���D��e�9���V;p`p$����9�#X�?&���c�Ũ��L�1�pօ���� ����y�/��#L�͛���&3�Ys#�� �v\�F�� ���xRr޽�{���̼`���è�=�vdj�/�����0�[�Ա DZ;�P[J�P���l7
k�޽��|Q4�,��a�͊`^f�K{z,���N�*��}�|ݖ�r{����O�~���믾m�?��<Hg��C4�b�*??6dj+v��v]��a��(n3P)���G�,�c�*��Q�r���4iP2_�J��iX��K��A��꭭�����6��������i�[;m�/��/� ���5'iĤ#ÿ�ӣUD��R��9��CC��§㜇0�`���wiS1���b��a{r��I��g���hb�u!65��čgX��ݭ�����WN	w��C~�����l:���ݤ��eV;������<�/��n�0�P�8O��ȫ	�[~2s	3���`p��_仺2����x�c2�cQ �k�v2{�?�w܏���x]�㷶����W�"�M"�7��m[ f��qL�*�Μ-2?q�(�-��+�S����L~ `��i�Z2Oi ��v�m��֑[=�d�䝢T9�Ht��s�4�%Ԁn��i�3c2��q�$��G�Y�ApR�{��5C}Y�	��%3J0O�9:N�͟�ڀ��µ��7����1�i̛)~O�.#�J���?�-��(�-����ԟ���������B����]��<��_9wݾ=Z��l*/��
K-�F�&���1xҶ�p'��.T��+LMZ {%Z��Y1Q%�
򆟵�ʓ�N��
2���}F����Z�6��P$�̓z�{�����u��Il;r ��]�t �ڥ�>�T�E.Hwe�t�ݶȆ�ޔ`��x���W[��z���i���7�����G�A�ˑ�@��U'^�I�V+RQH�S�K7obY\<�<\�O?������V)��=gP���"v�o�
đ������ �tS��3���|#ob��}vfo�6����Nw�c?ǭ���>�G��$ɨ게E��#&a�ON~�T�G#��O�^������U�4�Ϳ�P�0g����Hs�9x�n���S�q���J�!���۰G�����az��{ae�v���Q�=vWh}��1��mU�Ֆ��ɠ�؁w92�S����A���JV���y�����`�*�aϾ,[<ga��ŭ���-|�u�zgguO�Pv�}�ѵv�����ݷ��_({�ь�h㌉I��Pv�"A�� �P8c뽴ކ�p�@fk����%�b�E�<��*��D8�`�+�hp@U�ا�(��[�(�*��(����r�AC���ykK7��� Bp�D����s+E�ֻ��d@�!��D��QN��ā�wE�?y��}�1�I�`f�Ռ<��`c�=���b�i�#��8Y�e�X�^�0)�!y����3�t�6KY���FL'��Tn���j\X�
�Qn��2î���潬��C��A�zǉ���ŋ�ڙ3��ɓ'2��r%��8�i����.�Lg��@ KK�[ƪ(o���f{�l{޲� �e��g��,�)~�	��:���G�~��q{(7�zy:/x�`juI
�⪔[��#�R�7�޴յ���-��"�@���@�=��B(�!l�=��h>3�V)g�y�7�d0U���=�i?��`R�HC����.�3�����t��NS�^	[yX�RB��ɷ��;�����f
U�&��JI��*�ʕ?�k2�%�U*鯟�����?+���BYfx���ɸ���>K(o;C����D�FЎ�6��o:�����2��,�|��"�)e��C�
��Y?�Zm�:*e�0�fT�o�A'�
g�Ea~��~C��}f�/����e��3#ϡ���3����dFY��6ix��A��+.u�j���C_c=��v��qk[H��%<i�/�̱2ɋ�P?�{����>R;w3mg�SG�r[9*���C^���6�Uq~������n������k���]�@Z[{��C�Lj��h�r����mH�A4%�G�7�`+>��B>�p�h⅏��g徱�Am$If����ʏ�xR��Qqs����*:�����ʔ!�F�2���t��G��g���z�Ӭx֏�$�8��I.q�G�z�]ʭ|[y�H��l9�3������P����v���gQh�~Td�_�-���z��	KWCӷH'4�/�ٮ�IEa�����m;)	/��3q҆[�y%��M�<�h�ޯ�6��C�3������ߢ�~������ �t�����
X�?BO-��_������*��qB�=�}�=y�D;����Z� �l�Ax�4��
bm��Tij�������4*���v7���]�1o�|lhoFWb�y���J 
��x��p)чRE��;���(v+�W�=ޘ*�d��=K>�����1sI͌��;û�ɸ�au�r�]v�l>��[?�a�s��G�' w�� �?fn�\�:S����7��2�|;Aޅ�e2����o�����g��۷ڍW�勗���|#d�HV�k	��N�N�N��v���#���3k�[��g훯�o<i˯����V�_8)�UzD<�b��t��p��8q��?�]�t�]�z��3�4J�[$�*�cK��Z�\�E;tfD:m3xS�->��ڪ
����������v�޳���Mï�?��΃&��bw[Z�m
���L�Q(���oL%9�5��s��-�V�$���zX��geL�Ô����f�L���u�A�6yU~S"3ӝ�����|vez���; /嶔��,�:�p[����r��P�'���D��q��*�~t���[��3�C���ь�͵O�jpQ�l�z��I��%tS��@�ն@��������K���6�3�ݛ�̄n�/�t5I?ml������/��|���ݟ��-o��w���ڏ_:�N�8�N,��|���g�2�j�Ķ�&���q	���&���.���"�V�YM�:@�@���.�ā��� /.	ǐ/'�'g�kӷ�`�[gm��֣�Jۃ<%N�4�nl�dp�r���m
�%a,K�N8F ��Ƕ=�_9	OK��%LV>��w�R0Q�uO ^��Uf}
�KLcu����p=��]��t�
�I9���n�W@w���{|0#o�C�87��xʶ�u�{f~��}�)g~�w����܁���!����]n�>���F*_����u�߃�*���Z�ώ:Pe'�kf�v��x }��V��Ɔ��f��-'��׷2�= ]Eπ~}�����M���$P�&v����\"A�^�n�U��Y��OPn�������w�?j����x��Fk��"vi�4�nqoʭϥ؎���J��Q�q-��A���Rn��u�6�ҥ���"L[ qX������fn�ԩ���5gp}��!��J����J�u�J�&D��6`�[7�Z��%���t�K�w�,{���q�:]�Cn�mMO"�n�|7���5�}�f{l����+1Sc���#[�s�G%J�U����1\��?eW�9����^�<�gÍ�������nM�L8y��o�zv��Y�Tڅ��㏯�?�ɗ(��+W.��*_��ʀ��t0����n��\m��Sx�2�پ���ٟ��}��������2E�@��^p�0�݊��w3��p�ݺu�}����v�ʅv���(����ɏ��%�k�j/���p��ڕՍ(��|����헿��=}��2�"DƇXQneiL��8�:_$qi�g�@ˤ*�0��OI����{L���/�rƝ�+Ԭ�n�#��}�|�F�[ulq�#r��&��	��̥���*����Mz�hK��V9##��U(���	*D�Ȗr�x����n�r�L���*�~�c!J��|�,S��&qLU���� �B�7ʶ
�8���C0W!a�z�6Hq�����.H����7=���Wb��i&�2�>d�~U��^��]���a�ҥ�˞ڝ�ܫ~���������¹Qp�J�PFya����~�ߌFl���;��_^�l�z������J[A���v���p��7� �8Pv�l�����v�,��ٓ �������Ǐ�S'O���/�\Y�q[���ϔ���+]u��~M�Ӟ=_cp��=y�
<��&��S���4���o+��s��#G�N\I#���Z�aI0i[�Zޖ]����^��gt��y�5�
[��ߐeb:�{�:r����}�2�;�p�=~�����Gҭ��I6g��!�� $���3�z���9��~q'��c���<��q�l���	}�+��^u����b[:~~ZL�y����ڪ�.�v �*�����d�L����6л��7�ö�}�W��+t�Ul���d#㽆�Z�����`rV)����.�&���|W�%֤�ܩ�[�����������Oil/�(i *��h,r�8��[��m`�l=��=�^�! �'��:w���~@�֑�8�� �V���=��^�Gƣu�d����]W�6K�t��m�5mI�y�V�H�嵶�������ʨoj��u�!9�RoG3���:Æ�ښ�1x�_�y�^�����nl|�}�I�Ƀx����>|(��9�Br(�d�L��Y��7� ��]�[��<��L��/u-Ʉ�ktR���-��@H�,�Fr�	����|l"�_���O�?�������}�٭\	�'k��mm���<.^N� ^�N(?q�G��Tnwڷ�>l��?����_|��{��(zc3|Ҡ�x"٫�\�8�x�]�r�}���G?�?G���in�wB<\v�UX�ؽ1kc�JSy~�������_�x��������'�(2tp�7���N����4�)w�OF���&�#n�O�?�$�0��?�H�0OLq�F�J3�g�(�ñ��
_�	�D��Μ&��A733�h���1��<j`� ���KiƟ��� ��b�N�YVy�|���:���LK����f.io#�Ջ���:��G=w�l��C���t$�܊�*H�u�F:���-1�Ԫa(SV�R6~���;��[�'P�W0ߜ|�/@'T�͗:�~����@��3�)�����+F�Ig|�c����3���k�8��X��ڦnPn���u�R����'x�]�zn���j"�/\-�v K����-�ۇ�+�f��B�?R�����g���מ�Hn����<Lc��$������9��F�a�|�ݸy�}����WڅK��q���An)��_zM2�t���v"=!�2d��76޴ǏW�o~��}��p�۞�|����G�^�/���G��w�z�����c꽝��rf����S�V�"dd�ኯ̯��H|����7U��H�Y��#}�u0Y��o���>��Ƥ<�n��~Əs�'���Fy|6�k�?W�kFY����'G��o����׈y t+���T\�"�r�F%��Q�Ԣ��A,m��	����D�;w�t;s�T��yk�g��y+��d'��w)���67L��:8�D�u��3,˯�ۣG�ۓ�Os����:��N�"�����W��ۿ�֐������S=E��w]�e��n��`t	��z;���k��O_�\##�D��� �l)E!#ۃh�d?�EZ8���֖��0�J�3g��S(�� O�8��{r����֏0,��ks�-��~n[8:fw=t&�т�q �֕#�qVME��d'��<��(���Qbl�4�jt�a�t�ħs��ݏ��t��$U&v�&�� #\�����ˤ1 a�L+���П����@�yܰ���������<G�L�Mw��͟��褯��;.ip�<uN����u���O{߆=�S��[k4�7(���}~�V�v�\f\�l�
�7(�����q�� ?�+4�o	�l���f[~��=}���z���.���0R��rz�F�K�p��j@��x��>����+�ϷK��G�(x2kD'|�ߣസp�����.CE�r�_Gَ���Ez�b�=~���	��ۄ� �h\YD�aRS5����TךaZ�k}�:O��#��MU���;��ӛ�MM,��^��Xn��.��iƞ�A�gy��Mg��F��a~�e�q��(�+Ȫ(��(��
�xS�QV.�0��_:3�n��>E!<o�JiL6)�y�@����V%�J�>�U��Iߎ���;���N�W�O���k��R�M��Y4�O�����d�2�6���M������:��K��������G�4����� S/�C�,Ѧ.�?��{�����G�.u�=���}���� K'�?���}��b;y|�q�Ó\�&���~�HY[]���^�x��
��Ur�~�Cl�ʨ��oUJ\5�vg�.��~t�Z�y��������vڙ�cG���HG��}���jj�� w��;q�f�[�h����ݶ�,y�X�
�n9t��A���`�h5n���Jv%<+Vp�\~�)����?y��VW���fК�[��^c��Қ{���B��m����v`�2syɋ�iģ~�SJ|��>�]�!��7�ѯJ.�I�c�s�t��0��ۦ9WQ�?8�Cp�Ĥ���2��{������.���\j7�]jװ�]�@[8�"�|�8z���|�o�r��	���>�J����sgN�Y_��>�>��>�d$o�V����P�p�#��ܘ����}�J����r�;{������W�(�h׌�Bx"D�<̙���K[��O�?~�BM!�R�sgζ3(�'��S��p1
l}Y��X��e��ʯEF�F����:j��&w�aQ3��z5��FPDi�d
�HUc�'+6 �ء�t�Eˤ[?�^s� �����ܪb��f<���;��8hF��#0v^��v�^�@���^O{�5�'a|C�x�ã�;ŭ��3o=�BW��i¤��;�Pt��f�2���s<WA�pwg{K�r�]�t�}���v�ʫ㼑@��}gO�<k/PR�T��PEQ:����Ѭ�,#ԁ���4�_,���^�gO�"�c?��U��ڌ�\{�ܣ�X���ی��������Ξ=�.]<�N! ����eV���j��Xoۛ�m�T��b�TC��]��V��{�v�u{.e{��@��y��9��ˬNx�B�n)a�Vu3�@�Չ]�U�
)WM������{�GL�koXMw���+�t�e]�{I�)L)���t+Yj�_�<�}Ј�	�k�t�+�;_�B���l���Cu,�/�>r����%N͠����hS+*��<��;��Jfn��'�m]���
��L98���I/oE��gX廫�I^ΐ���l��M�(���W��,5f1��<H�"�#@����}�$d"���w7#��T��J��8�*�ʭ�:O�à���q��ȋ���m�6�~�r�f_�V�V��j�7��0����~m�=u�m�� n��z��={�,������˶���w�ؚ��W�l��k2�>����è(��Q�ďE���;��H9��6 �H�ݪՂ�M���٭�_ڄ�C�J*ke�����������#ɫ���Y>q�0� ^-�"K��h)���s�n)%�=m�^�ޕ_�@��H��C��H_�>�)�}���K�l[sf.���0�����n�M_:~eww�|t�O����u������d�C�3�����˒�L���O�6�� �[?�Rl�9S{�]�p:�ҵk�]m7�]���.�Ԟ;s������-�S!�NP:�H��$�:�1��s�����=�`�A��A��(���nz�+= k�g���ȃ��,��Pi�ڑ��c�T�^l#�Ϟn�������Rnm�F6B����K�6X�:�-��1:�#9��6�V�S�g@��������J���`rgmWd}W�u�o�ܖ�Y�91'�֎C\�A(w��7�C��-�����Y���`:��k�>������9��f�����W���f�y�_Q:��ٟ����ߐ֞��S:��F���[L��7��<W�F�GF-d�[���l�d02ѿ�
:�٠�1�_�=�خ\>�>�u��{6��������oOPT��������ڲ��R�������`_}���XA�]G�ݡ�PX���HϜ9���ji��Ш�f,�>N�>�8��H��}N�����Q�W��VP�7ȿ[G�����>�/P��>��o��Q�@-������:P���imM�V��J��A9g�ԇ� �^����^�����k�K�7DR�'�@����<S�H�7��~ڿ0�����G�Y8�C��{<��R��mn�pI��U������ํ!�<�+��A75n]i�LWn}��	�RZ
m��U[�K<���r��*I���<rȰ�� ��\�J� �$m�h�O�R	#n$j���Oz������=&I%���!c@) �V��V�
&��̙Sώ���A�͛�i�'鷬����U}��	J�K��M��6��.��L���L���V��͍�L�~��I�ϟ���{�P��nCO�;��������+L��C=5���*)"ʥu�
�����<�Lj�<0���R��f�Ú ��oȟ����j{��y{��q�ʭ���J�����������F�yɻN�}wU)'�Q�m3�!�#}K��C3� 3�<���6��!c@��oG��_!�ʹla�?R� i+a)��^�n|V�Pϰ����n�k�2���������π�|�qXoc��ɖ#���%����GQh�\������^G��~�r�t�|;떄~^J�KEٺ*�yѱ�G�˒�q�!�ț��z���'O�؞<�}���$Zf������<
�&�-P��A�ak�G�ɥ�s{�T;�W��Rn���QɈ`:��7� s�W���񫅻�����S�g ����ԋ(.w���cκ��.-�wgi�V��|�$��L�>0�3���l����J��qK8W\�l��42�n�(x(��/�J$
=nKH��k��~S���at��4��_ʔ������`�}x��� 
&��F����[�t��1�j$^�|i��Þ���a��[RW��b��dR�+,�4����w���~�����ꕋ�[7P<ϐ���T��s����?�%��Q�q���4�����d�XY^�ҹ����_��Ф�o�/D8�G�TyK�����p��u"K��/��p��gy���.뭓��s֧��D�>|�/��|��u?�+�x��A��~�w�.x�V��H6�j��ǯ�Cgn餲�^���=����(%���FR�E��ofF���ה���ă��}��3mU�❽x�=;�@�@����H2a�1%��,Ċ��ܡN4c�{O���?y�=�ʳ���O�0�ZH��ȩ!�ͩ#bz"���cXq1�(�(�5��K�qf�6'�I��zW��E���o���ܒ�aǾ��K��B%�0���O����g�:ό�������Ƭ�q(>*�a���Rn�}u��E?��_8I��ݺu��;w��<���
���o�o�����0+>��?�0����䭶��֞3 }��q��n���oQ�#O^������V&�*�,��Z�4:(�w�5uU���I�w����^�������F~���׵�����
����/��3����S�G�!��ř��V��A��-��uc(�$���d�!d�	�r9x��C��9s��:�@���䟃��tC�ue�/���e/�=�i���~z�	�1_xp�?h?ח|����+����ۣi����4�୮���NP:D��f�(#ߕy{�tY�1�����&��aWN�U��r���q���j�Ph�_�_k7n^˳g@.�?�N�<]��²زˌ63@?M���m@���ʹRv����#�p{qѾ�h�خ18�0�+�ʲ]����ҕ�R�C�N�;t�T]uѽ����_��?� ��6xZ;	����(�C�U��V�FN�[[�4�'5K�U#��R�l'@�;Z��?@)�C����&�Z�����׸G�5��%M��Ť6��tv����fWs�~@���>�>o
�y���Γ�{x�>e�{�1���9�w��V��N����1��{�q��?����FA�kLe%��V{h�yp�ky͌gGQ���v�������Nτ/�����v��{��|����Sn�?���*����s���e�r��Q����2*���9v.���[!�����R���W] ��r��
�#a���-�[VV��l'����I	���ѓl���a�s܏{Xs�XۦS}��N��+�`�ܢ���!��m�E���1����D�͔�0�=L���Y���`��C�)�8�\< �zN��%���Is��x�}M�n�)�8 +�u�lR�`��H����V���َ(�vꁥO��)��IzϗʹU"���%�O���3�����M��|��Ŷ��L��ɚ�ݫ('�lK��/���,whO����~Ɍ4R�Q���<b�~�?�{���ُ�D�9��� ˬb벺�����v���v�څ(�*j��/_�j���7�o�{�U���Я-1H>��Ӟ��?Y_�@�]&���Oۋ���c��J�!�	�E��V[�o�*�E�G�]Zj��s��W9��v��-
N>����~,����L����[���V�r���mY��v&�;M�?�����=|�V�֠i"C�/ _�E�v���v���ͫ�����"2�������δ3(JI_�UQ|m�����3�J�l]����>ui_��,�?d���>dL{@2�nØ'����cVrK��"Ws't
�K����fz��O�.�f�|����ΠL����������Z�����ƕ@GPxO�X�:K���^�2�L핫���K5��Y�1S[[��,��׀Y�����+����.�~��U�㜨Q����b�[d�<m"E��~:�W�<�A詮jD���{����2�������K Oy�G#3�*����a��E�u�������T��f��5s�m	cú����ܡ��,"M�;1%D����SDʻ�D��TT��x�����C¥+��-e���m%��4��Qp'��?y���c���7`�����|��g@lG�ۻ�u3�(�x�f$'M|H:��g�͘��<���c��LKZ�	Ae���Cb[��W����cD1�<���3�ʭ{�Οw��<��wi�Y�gO��x��޹K��v��0�E�|�օM��/r�}��Q:7ğ���4������3�'y<�;����Ut�Pwf�CcW._��Jq���q��x[��x��}�\-�*\N�:�Ν�������vN�>{��={�,4=w�"x�i'NϬѓ��(�����g(�t\�Y�Тٌy��֕OQ~BS���:&���L�e���{a���=A����7�V|5be}g��ǌ�~g�����soM-O��+�E��e�S�l2*��C��q,�e����B"�{8^���m�_m�p�9�:s(��	�eH�����DAhMؑ�!}����LV)��j,��G슗�{~&W��Ch�������k��5������*���j�VE�����WGh������-���r��~��۽����b?v��r�*m����'�X:Pv��=�[[^�K�w�.m�qVr�>r�Oһ��P;I�gr�gYQ�|Μ4;0v���_t �$}^�(���$s��˿�9����%ɏ$���EA8�\�m��Vw���5@~��Y�WyVF�(p�|�|����G_~�~����/n��o_C����>��J����O��(P�/]F�y��1pE3w�9
.|�^��Ͳ?Y=���g�T�1ư��~�1��U��z1^�'� l&��]]E=#+2�=�g��m:�np��� s&N�������
����0]V���-)��o!.^gP�`�㏮�/>�����f�I�������0�	W�)�J����6*��.�Gz㟬�H�n��S�8��~<k��<��|iKb�7	Tj=3&��_���Y/�Vb�	G/
��: S������,��ښ����X��=�����-�\�[��3�O�R����vP���؎0�EP�����z=�S�
}�V�3���h���cj@u�Ť�Ԩ��$xeŴ5�Qe}�d6Z���N:�gM��G�83��<L�n�¿Ew��üG	;��	�4?�֔��yf|�G��biU�r
���mr���_&.�v�C=�Z�ø�.T��4ع��iq�J�Cǯb��4f��ɟ��!��n޸�e3��wP�>G�?m�>L�s����>8��6����m}u-ʭJ���i[I:S�rO��p�����n��S�*�n9�p�I ﴍ��:��O���=҅�?�]����s�η�����~��Kg�^e���~	���s�xa�(��i[^ބF6`	G=0�yCH��C�<�ό��&�������y��)���� $@ۿT��̿�53��Gt�<�%N:��<g�w�͛Q�2򔲢�f&�1vd��T�q Y���a�y��[;t�ϝt�.*�1s;E'9�%8t �PJ�լ-���Q�O�H���#��C6ߑg/G���AZDØ/���zY���t�S�ʣh�!��s���<�����tz�L�p����]����|�l�z�2�H��~��}��w�5gΞE�����)
}�rt����W�bk��Y�J�n[R�uF6W�qe� 2�0*�����"�gUp]!����>?�<B�(O�*�l9�����`�B���X��/�zߨ
����˗�7'3��v���^e[�����*�6ჷ�0\8��z����V�&���Kg�r�jS&��wNt9�� �}�90N���m?b�Y�G��4U��z�3��`�f���)�x�]Sq����1#�����W����@z����X�=�V�#̈\��wi#�`�-U�TQ����Ү���Q��X/���>��ʝ�EY��`�zc�$�}|�Z�����!J-|�Ƕ���C��-9�wdu���y�SѦK��E���0U`�˟�sF��zXxUP����V��N�#Ok{H�QO�����\ ����w��秫+��\wc}#��ܢ${���l��&��{mh`g!�U�8�e��(6��m	0z��ip���� ܩ��Τ�W���A���L)�S�Q3���|6�3ߙ���Tn�y��u�ت�"�0��r��n��9g������n=Δ~9����M��E�TG�{چ�|l��������,�{�b�����N2�ň�?>� �@�$9F^����n�<cRr��l(��%�{�����8z��������O?�r��0����f��������:�j�+�
���a]��	a�xJ��c� ��D�u@?X�8��4���A��>�tJ��w����5C�>`:�3�-������u�md��ߐw����Ip�̭��hw�>i�w[B1�0B.DL�r�~����p���`5Ͻ��k��&��ca�-�	�r�x�_�]���ϰ��/ςQG擌bF�2�6����^wyi"l{:��FZ�{�E^� ���P�ihj��L/���3l%�T�K�vcv#�iG	!��T�f�d2w��3��#|�Ē�6��^U�
;�$���f��d�H&��t0.q�|�_���J����z7��/�Tx�G�T�8���f�|Q��4�B>�B� ك6��6�����=́��gζ7��Ͽ��0�鸶��^ g�am�%9�$��u$=�*y@M��Zi9��-���v%��3�'�!��RpUlK�=I�3�㲿�4��b�
�3�nOp��[-�{O�:y�!oy��+��hg���៍��v�m	(�N,#�4�@�	�r�|��OPlo�ПG��̣��Ұv��u��ۤ��r���uU�8E�}��֝I+CH��<�U�Վ�I�}ؤF��{L�ϥc>��<��V����D7
�}�^����;z#�K�q���n�QN�y�j�$�q���S�m�SZ���;�V�ր�jy^~�y�J������^�ϝA?�a?�p(�ڕY�D<$�8Y���x��o��l�Q����I��:��1�/��EN ��"��u/O{��L�u���&�9빘#�te��	<bUH%�«��u	�H���
KcĨ�y+��[o<��N��,㑮�gf|.ȟĚ����_8Z1��q�0��
�6�5�P�νC�m�-A�<���	��_!�a��O�g����<��}�3Gɞ���A���b��C���T�4i���~T &�ͥ�|����π4$1������[a�*Kf�p���2\4�ߜ�Z����Qg9N8�� L�oÍ0�#I-�vnOpf�=r�� G���u����R�=�;�Ess+�@Zb�Q4�Q>e�M~���su�Ի�l?
���E`z�����;rěB�Vφ���#)�����w�vBa�A��f�%-$X׳f���Pf>�2���R'ZA�/�q/4�`�R�fV�����Љ��S	�J����l�,�g�K�!̇�V�pӇ ;:�i���Z�$iN駃��n�=P��M�,�	8s�w۞���t��4XiB�Op��gx;W3\��Y��Lo��c���T�`��� 莭HMY;�c����i���/����][ނ&��=�2���$
ㅋ��C�tF�a}o�����+m{c�4^�c����-	�ݻ��h;u�p;y�P�3'��=�Ο>�.�Y
�G�={je�aܶp�4�_M��Ջ����Prϐ�b���4����lyonC�Ԡy�=�t�72���S���)���>+���Ϟ=��y��ӗ����|�}�կ�m�����po����ewwEz1�k=��2�l���F�����M�����՘%�Ly�L�w��%
��4]�^k������N=��1@z��I=x��π�����d0/��T�x��Va�}_h����o�#<@��.\8���p1��@I��U��G~�|�_�������d؂�.�R���K�A�
�k��g�[��+em̸�%�X��[7���>��>�}�]�F;{2��Rޅ�i��)Y9��.��E&�X=�	�g�k?l u���e�L*b��s��cc���AUp1�5�B�30���$`E���fcא�^��y���,Y�������'#�5�Aa�C$�>��?!ӓ�P�o�2�������`��8g�;��w�?�o���X~�W��)-����
����7�u��+�H� ����d�i�Ζb��Tp-��^�l	8�GE�&C<�KN���F<��(*�
x�YۂRZ��q$���ٶ�fg��mu5��'���<%�K��og�\����(�z3��ͮ��x)d,��
;��eV!���LD�=Y�}F�+sb�z��qz|S<����{a���'�wŚLe3�����xt�pe*��&���Q�C���	��M�g��"W�k���{��'�Zų��l�SF>%mӲ~s�BY�Bj�{�J�#�.����ƫt��+��!Ql�ð�
m)����_#�`��j����ƈ�M]{���s	����s(
�OeIb���]�Ͷ�����W��b	��a{��Y�Ey�1��G�Jɡ�����}���.��7����v;��5a�] ����WOIWy�b���e[A�u�Ǚf;b�͋(���W�)A�?7.Ǆ?��O�v� �#��k=������r��Ͼj�����������q�;�ﵿ�w�������Q�{�����?��v�{�+��B��������.�%�ɋ����\�XF�y��/dL���^�O:e���c��)��8t��k�֑�k�kt���~���7����E�����l�^;�EW��t��m��o(.4�Ӣt��p7�ʪ״���w5��R����|�I��q���]��:4��}���KeJ�4�峌�9p��i�b��Gy�--*��||#J�B��T�-�P�Uz�-[\*I�2����t�fB�I��~�i��8���El��R!T��-�E�6v�pgV��]>h��33އ[V�D���^
l-g�eV7�R�8=E'{�it�I��8O���$��93��߿�!��p$�����}���!����Pl�Y����ܓH����E-n3�2�/4Y��0�?G�Si��]�_�r*���/���)�N�u���,�P�6�l:2���;ʢBGP�*�e�nTjO��+JCV��
B�4tӫ4�Т�]
�
Ie}�aF"���R��g�G��m�v^N)y��<�D�n[�*s��d�v>|����?o�p f��t�)y���e��F�v�Ln��&�z����K��5�n�P`+�k��+���\~�u��{�!���$ʰ8�꬞S��\�n�
"����:�ԽY���oOp��ٙ���w���x/�<��h���q�@wi{>�9�烬���'dz��x'��������_gr��R�[���ζˈ
��o�G��]p���I��54�Z�!�CN� �9�̢��I]���02�+��s�x./g"�Ώ��l������k� �����z}[n����"3�k�(�E>�w*{_S�����������w��������_����/ڟ�ٯڟ��W�׿��ݿ��-/����Ň���m���� J.�W�:�>ƞ����/hL�(�YZ!0�]ꋐVh�?t`��~����x��t���8�.�?�y��?��Ξ>V[KN�/-��O�*ǯU�hd�h�{�h���̗?L���G���~X=�3 �����(���v�B}��$-�e(p���y�W�4�%�U��1)�@\���2"�f��Κ
g^�n�hc�u�y�R�<Wh^` �b�s�a�����|v��ykۯ5����#��oI���;���H`|�/�+�0�i��9!l�@��3��J��T�y(��A*���%�T򅌾�Yf�A��D�_)�)����R &��!����e���0}S�
���o5�q>�}������ �%e@y6�;����D���i�̼/ڠK)��9���7��<��[�ØC�U�f���졊����;�����S�f= v�o�π�k����FfD�{��V'��?q)����0Q،�bt��yԶ�<�U���y��ʃ��`�XI�z&�|YJ��J�6c$��s�M0U*Pd>�_
�4e�n{���Q\��߉o��@�7�gf�;��K�@��^��Ѯ���o��3��I�Ң�T�vPv���:�\C�7V3]�/�G�U��+<�
�����4��h+)�|H�w���h�a��s�Pq�WZ3�-<v��p�ߙ^g���Jb�? x�w��we�����2�����7)��a+S���&��_sf�(��nK�+����@�@���#n�����j���FX�B����������K�ҳgTPj�]�*�n�s���j�fȌ���V�uF]�5X�ڴ�Nm����C�G�c�����y ���W���g���W���Z��wu��)�����u=�ܖ*R���*:P,|��[S!������ݽ6��=�:����~�0O��%��S��s�O.��?�Ҿ��Z��g���g���۟\��B�p�$J0�����lQn��K�ͼ���c	>>��=t�g�o>��5��(��9����CL�������5鎙�Rt�Md����#X�'ZG��_���@��f��SB%^���G�+�L��6К��r��{o�{��on�s`(��)-�cz>��Υ3g�d���aD.�ʽ|(�.���ft��~lGG����B��2���f�;��3kg�Źfgk���Q���4�B �)�,�
�e�w�����y�>ü?)��a��a3����8�F�1:q���������fbv��3ǘŤ��W�ށg���WA��䦮��ޕ���2s�,c[��QZ�38�bˠ�<P{{��A���������K�q���;e�>{���د�V-����f[�R�K�{�R�7��}�oYM"-J��d�|ҭ�.F��p��a��ӗ2�#f�1{���c��q�r��\�yϘ��fV�n�v�P44����� �p��C��d𵾨 ���F�_��ī�����Y�4��[R#|�uI�U.;�/���<z"��f?�����/��nm7Ȭ�y�݀�+���+���Yt�����=�ߎ�0��X�ݞ�jG�B���օu����@;��qh��/O�˄ȋ��c<��I�7�@���6�5h��j�Ԡ'�ecվ\��/?���F�ɇ8�$g;�u�C���خ\X�*������qn4���Š��a�����S��EE۔vm3�c����S�T���A>��CSi�B8~�?��5��[4v��*����%��3��Pj��?����?���?����|�ɏo�/�Q���ܽ�uoG�lQa����T��Ky�[��4��A>�U'#�����[gm��û�?	'��RK��N�Vx�����`Ն��q����ϧ!Lf*����"�������&�$x�Rӭ-ꤰt�0=l�L����skݍҎ(<��H���9����^:�F*��G	�Ag��"�~4����ļ%��������e&"�����e�1;;\�R����)�3x�O�]��-�](��+��)(xW�" ^E�@�8���1�y�2J���2o��H[� ����w��o����]���֗w�����W�6{���U̿W�'np�C��C25�O]�F��X�֬.�^u��1xAE� �� }4i�a|Q����i[[m�OWf�c��ՠ���u����8xR�_ !"���b�~ّ)�*��L�Qv���K%��ޓ�^�7>:��L�E|�W�' ���X)�-0�=�[�3W�;���ںWۓ��[�m�;38m.���}�>dHdC_&�h��!��0ݐ�^����h}�����O@�6��:BT��?�GL.���[�4�f=�0�,�R����^�-e���i��P����I���?�G����T��m�(�V��0���ȯ{MP����?Ŧ�S �{�S�ӡ����p!"�����י�jrȗ�P</�*7��v����+�v���Z2^J���7=ۭUV
��~�?u�Z����r�m)]ڍ�a�$�e��/n2����L���������v��b�r�J�v�f;�r;q�,yz��[����o�w���Z���|6�𮃾���c�'�f�g��}~¬�L0�$�� �:�7#xHˏjx�����j?���ڟ����������_�g����/������?�Q����v�ʅv����3�哐�4Qnmc��C�U	��ͽǍ��a�t�!�Ν�K��B�I�b�*�����EdɌ&�L����}�Et3^�#o��>/����8 ���ۼ�N�q&o9zĉW�ݛ���ǴG���&	m�����(V64p�᲋���BS�"���Xs�P)�G���J��2	��t��g�1�օ��9Sb����fg�j_�#\��f|�s��׭*P�iM+e42m�m�� x�ΠE�=�J�1I�MӿJ�}0^�� ��L駪g�:L�����p����פ�M��q�{`dS�1`>�P�|�?���[�U�358���IL�`4�f���}��thPo�
A�Ѹ����D\f�;N)p�m���E��j+me��l�(�[4��ħ�i�o��7ﯡ��o�x��!8�T��m�Mԭ�g���^V�/<kG��,��E�C#~�����,S:%���έ�P���=R���,�2��_0���Tn�a��Э�>9�?�!��O}Y��Rd�B�f����z.� �،pS�i���.����߿R�����)��78���[�^qr�"u-���)�-�K*<��Z����M�&?q7j"7���
5�T���K�#�2I���ԗmS���*ۤ�%�^���3���֔����1��7L|��'"�����S$�Vi�=m�|�>��e�IK��"+^3�v�kB����QhAG�����ڕ�d���,M�g��5no�H����"+ԪM�5�y[+JΖZ�BRk���W剐��)�O�m�P9���e�����a�;}�t;w�\�3�Ņ<�N��V�s���豥@{�r-_�|��E��(?}�&>bUy�W/ǐC���c��p�`�� ����i'y�:���~�n^n�}r#��M���Ջg��g�5��ϷW/n]��>�u�}�W�._$����_r��&���Yr{�	bez==D�:�A@#���n!��cQjݎ�2��U�J'M3i�C7��\���)�
�߇���L�)9�{������'�2�M
~���q�4���A�ˢ����1#c���w�!Hd���f�����z%�Q�)qG39����Za0�#O;VƱ!�0�)�/����!3������cK4��#�Z&t��}�G���@by @y<��R�]�B�C�;�n��0@��5���
���V�h*zf��N�� �O��r���2�RO@�EB���3<�'�:�©���	���:M�*��G9���|�߄j0�y����c�č��������[g�h�F��p_�3Q�oz֏�JH�Q8���W+����:J�n��d��v�ސ�mrŋ��ց���*����.T|�C�m��vV�:�)�c�cQ�U��	�����o�Wk�m�o�o83�%W����v~U�vVMQ/5�EY&?gQ��uY�û��d>� Ӻ��҂�C�"&�{%t����Sc8�����_�U0��P~�L�f0��Y{�8T�2�p�_��Rj���a��F� �����!1�u��0���]X�Hx�#t�	"P8�2V0�ӝ��1\�?���|�P�I��f[	:��C�e��Lh��_G��i;�2�&��̝��#�F��v� h
qmF{�v@�E���c���<̻:��K��w�y;q*:���	�WL0��Sx�,
|��!&EG�b�P'E��9f�&�����l�Fbڡ�}��y�!�(Y&�Hى�#�G �s��_#hۯ���ey�*9���\D	�P
�v�d�29pp�x;xl��c�푅��l�$�M�t���tVQ����n����K�G>m!��\^�:�_T޵��o#�v��֝�v��Mېrhum��p�ݻ��=�F�o�¡��ҭk�I;[#����_o�����g������'O���թ��@��x;�?rK�݈��Qwc��i(F��u�g�]S�Re�=�ׯ_n_~�I�񗷣�^D�=�r�zs���&��כ��	�C�'ڍ+�g�j������Y���\l�����T?�o
�fVdE��#��*�(�$�5;?��T�_+{�~��'�x���Q�}V;���to��V�|��p#���M�4�J�U<�F[JW0md=�������'����d����;._���ӫ��><����~�M�͒#hedA"�������:���A�Mg?��v�FtA*G��*�u�Ǝ&�?
�	�����^�/�0x_�ak� w�S0�ٜԎd �+C���oc��
"��_	�yP��f<�"���1�ۚ��~Sn�䁓��)�`����7�n�Ѓ`�����w�$��(���"��s�F�O!�g ��ʝ�3���e�H�4��A�D��v��yβQ�%�GU���|����y�ͧ�^-���/���T��� ��h*��t���������+��2�ndT���F{���u{=a��$�>��aUjK��ߴ�� M���Fۤ��"��tT*��G�@7i�E=�lJ��=�\��#��7SB�1��z��6�)桛�{iO�]PA��A|t��T0�x��t<��{L�Tm�n�W��=8%8�GyF�I1��N���(���Jn��4!�s�$�w>}e�~	�bM}t|�r��c��g9�w�%�rY<e�r�ˁ�m�w ��$4�ߤ<�Ƃm*�swC�N凿&���]3�-�~��&X��¥��<�d�r�%$��w�az���}S����~�Ұ1�(���:P9��Q��p��=v�[Bi���Cȕ7j����&㭶A�-�Ҧ<`��ma�[o�9�ϻ��
��>��Jk��##6x.������ۍ��@�y���]Ã���)�n/��r$u�o�e��V7�u��
�,��76��>x�=}��� ۔���GX�(�m}�KZ9���/>|���}�r��={�<[y�u�`�j2Vn��I��50/�~O���>�j'Ld�ʞQ�=x��Y���{�|�|�l>d�D�z��͖J�F�u��:J��.u~������v�B�u�j�~�2ʭ�P�-�.l�D2���̷�n:�������zʗ5O�h����S�i9X�C���=?i3����3��޶/q��������|�w�W�r]=�jŰ���h~5��8s댴q��J`]��PƁ�A3H��"�:�L2-�0J�q��\/i}�B�?h�B=�1r����<�Lʝ�9�o*o���&n
3���y_2�3#��;{��5��w3���<�>Ͻ~Ȍz���������ƆY��
,;�ޱ���44�S|H���賲;
g�of�d;����u��٪�c!o�Y�l�*BJoҠÉ�KFJ�$w A��^�Zi���h���(�tnp�[���D�L����'����v���� x�P��%�K�_�{������{Ծ��}����u�A��~���hO���Zo�^����?!��(��tl������p�3��
�R����ݸ�G�� -��d�^�����hY��K�*0?h��4�+����&�����K�|`8�+(��n�aP�P�j�#u�@ɺ'e[.�:���?������Y8Zn�ә����Ar�e�I���>	=�(��Q)��rn����dt�,&�8���E�62�}X��OϘd�$�Ồ=�駜6\g�=`�c���y�W��7�P#=�?z���vc�D���ɧ/��3��s/��w P��� ���A�� ���ӹf�������~�t7+)��t�x;y�T;��KKt��PDwஶ'/_�^^�@�U!U�}�V7^��6��l�o����r}�=_�iO_m1��l�5������C�g/(#��!��w����ډ��۩�(R(9(ܮ@Z�����L蕁�
���+5 ��Q#~2ׯ<>|�xО>}��d��]^��gOk�[.v��:�}ه(�w�������=z����[�m���)GCA��{yZ}�v3` �a��!u.�h;�<���b�r{�J��lo��փ��v�L�a�����mcm��l�_��c�ڙ3K�̻�Μ=Ezn�p����������#��qӋ��Z�*'��������\��>�F��� Z�Dw��N�:�߈�0C���0�?�se�<O�[�+��^q&X~��|	��l��
5 ��b�dGe 8]���[���X��Y*�^���	V��;������$GF�<�/��~g���9�o�pxǣ���wPf0�~��&A����3J���۱���a���iO;n�Z�4K!��Ħ�[��#�}6D
��0VhF+����啕u���%�ɳeX��.b�=p(�v.�ml:˻eV%T���y{�d�x�=|���{�ݹ��}�����_��.�}���������7ڝ��+��/Unג�}ۇ(��p_�p6E����=F���ɑ��8�,�++�Qr�sk��N	�H�h�� �D����6�?�|�y�9��k�wa�y���Dȫ���U8O��rg'���À��9vW~����Еޮ �"�HY���@�܊�<
����\U!L��/+5s;�n�h�W3���!� H%h���v�D(�:D��^��Ҟ��!#!�"fo>U�hf�퇞s[�WO���KA`'e�+;�m%q��e}�涘?rt�D;y�L;~�t;|�X�,=gP}�Q���{̠����>~�<y���e�,�{�V�݇��}�<Yk��m��n�Т`�ڎz��e��+��]-�r{t�-?��@K%]9��,���mkR�T��Yie)3�/-�.��Xul��*R�9+8�~�Ѿ+��S����m�4^ߛ��cS0?�ZwL�c�f|���4�Ӳ���y]�Nh�Ok�Ν���gET`\R��=��2{0�����kE~�m![TlO�<�푶�1�Rz����?�>o*��O9B|ie(���z3�w��0!y%ޞ�T�i�[���4��]���~Z��[���odYK?H�˽��i���D�#�è�~@ږ��嵂�婚%�;����3xh��.h����ϛ��O��ެGOֵ� %:� ���%�>66ַ4�]����ݎ�J��s4L�4Pi͸m��m�`��2�2�eh�yӽ|�/��%^�Cd��2��E�Cw�e��k��=z�?yіW��q�ߑ4
�k:�-��m��/������w۝;tH����Oׁ:�U��o�_��n��?����}����ߵ���o���]��o�o�{���7�����Z@��!8x	�S�ەUgR���"e���{$�С� .���	����=ᶻP��pV�N�� �������K9YΙ��ؔ�����'�)3�>`"H�;LfȒљ�:�͏��%tE�JvL3�sp�?�YNۧ����0�Uz=i�>�Llh^2�f�2TP2R�!8��v�!�)L�R@�<E	�Pg�l�)ۗvpƯ�߉cZSzs0����~�������y�M?�|j6i@���?�F��Ky ���������P�MU�ݥ>׶�e]�v�u�R���-\8Ԏ�Xl�Ν.�c�O���������U�G?�u����m���^��Σ���-�|������o�����������{Ѿ����a@���6����[�~����W�\M�F�>z�]<%�ܑ{�o���7�:J�e��+�>��;ی���V@j0}��
���瀳�!���7(�����W���Jۂ.*xD�R�GΞ9�f�N���%��9��E�Mƣ-�\U7�D��V1G)}�����	�;�1�Ν�}�Kǽ_~?9(~��JN�w�l޻������=�n�e���_ci��R��j�gE7M�!�;�����ٯg[��͈�������s�ު��*�
[��rSe? X���x�B��d� ����"�#���[y3o�i�D�w��#�~�c������{�5~��f7�c�c�5�\�#���8
�2��0����'����v �G�|���q�.�Ү�X}5�#�����.Q)�\i�|j;hz'����EU��6��Z �A`R��@�a�4��@���k'8���Jى_� � ԃ�@t� ��s��1I���F��ɟ;�T��Tb�#+�t�X�39Yu��@��?&W	~ �xȤ}�����Jy��&�U+�+oQ2��x�J��/;;�e{{�[66���:�_�7e��l��Y�)/5)={�V�H���ɲWq�H�}��穔�/W�j���[������ol��o۸�����?�5!I�=8dši�WV������hΔ�Т?�@�p*�YnU�e7���x�؅t����_�eZ٥�:C�0��/Y�UR���zb%O�݈]�f��) %%�ˬ�1VXq�c^�kĝq�uM��ɸ4�~L@L�񈍶^Q��q\Ҵ�L�ɏ6&��+%��ղ��e%R'��vT�B�!���t�uҢ*	-[�IE���v�H���ڴ������o#?�ȉڛz����#��&:v;������G��8��u�]F�G���|Y�~�,^�^&g��M���֬���1�n���\//�H�]�*��l���a~�|]��0Vf�ؾ����qY]?*+�O��G�����������[?b�b{�����W���-S/5�	�,��س�T��mO�wʇ�pU����MMM����͛7���#��k<�Ѻ��c�2G�i\a��R2;3�c���!�u)��Vziӱ�ɹ�<!V��n֟�x!�_��l��zdD�E��Lt���V�p��꼹�.OjXET��-N���rE7�%�@��EE�G��X[�O
�m�l�)�ԡ�P�,v����1�;+�q�Mb�e3y6��m���������@�Q7m�tl�����˺`�1���c)����) �fލ�!n��a��� k&0d�i&t�>Y𵤸��k������d_�jr�I�qw�Ԭ����H��x�Ǽ^��X��Q��o�V��w�L��x��!��n�;z)g��zu�؏����n�:�3� ��QluAI`�$��f���������o���|��w嫯�)�~���|�J��&�����N΋�rt\�X���-��`�Ԥ#%\Y��D�NY�һ�	hee��]��۝ݣ�'����T|Nʮ&�m)�[�����vٖB}��ߗݽ+���~��]^YV�}M���ƪ5O�<N�`U��-}��*a����rJ��{�j�Ox���mD��bi��cM�9^]��ɹ��aVbۤ��,��P�r����"�iO$�b��]�Cx��z��������ċ䭮ǖ��o���@C6��i�9�=!�3�*��l#� ���,��);��4ۮ���&^�(���B��_	(ٸ���f�<�?�� W;�ž��V[cZd���)+�j[�s�dw}p�ŧg/{���1�j|8{WΔ�ڋ
g�.,͕[wn�{�?)7o�/SӋ�7��~,%T7�Rf_�ٷ�%V}}u�[���bG�}�v���c�<I:��-M�ߐҺn����Bq�����7��~^���i����o�����_]��������1�{�ؿ){��RFU6.� �b<����BD�RF�???W�߻W>yx�ܺ�P�f�T&RP��)��253^�g'��O��bڨW<?yx����{�O�۷n���q���r��_��#��8��t�.���J��Wy99���<1�؛�VV���ځ�i�[ʋ�YP(�'ʄn �Q�=���m#z�~?��'*[��.��������8<2��V^�/�Q�P뗌#j��bG���놶9bl�}�Έ�e6�~��|Z�4^��,�(s�0�L�4:tawa%��b�\@ŏ�s&�:8[L��6,�R�F^��� a��n$��T����I��gK�E��W�����i5�A�!la���������`(�401��]M?�I��ip'�c0�Ѳz�)�J�����V0:� ��c����~e2�H�\)O4|����o5�3���W���7�e	��~px"e�\J�l����C��ֱ�v�^"/�]�d�?��j���������x[�R���o��6V�����@�,��NY]�(ox���Jy��uy,�g���v����S�n�o�[����� (g��_o=�$� ��c�����P+���~Q�NN�J�>�y�:&ϢQ��1)�$L_D�i��_Ea���h@�}*� �Jf��%*����*+�(�PH#+�:�@�ﭥ߰
T�>@H�o^�/g��i� cY��G/� ��Gƃ�1.@�S�������@��9�v�i��SՉ�f��$��rմQb}�#7O�y�B{��?+�lQx_��5>l���s�ѧ�^�g/��Q�@Z_�ݱ�ӳK�������M17���ek�l�/�{��=�T�����e�-3��w���U���])��y~���u�ek�!�̘����巿�}����m�'Rj�ɟ�����Z���ʓ'O˪ƶ��#�'J[U����2mQ��eX�XʊU3�s.--���+�|�qssM7������O�;wn�7�� _�xxT�T�gezj�\�:Wn�KS��wJ��OB
Z5�~Ѷ@T�+�z�v�^�d�(���&��j"�5�iح*��4^D��������)W��>,3�Z8~���<h��ю���̣_-vƀ@�cܐ��EQ�/Q2�!�<�_?/����4��5�1v��f����Q�T������  ��IDAT�������Hw����1!d4���K��QĈ&�0�h	�ȏ�k�úk�]��AP�!�9�H(�XYYz&�M,]�	O�P�L|F�X����Q�t���s Q`vvP2x#]w���r�;G�ҁLѩʈ�Ҧ��>���F6{ָQ�c�_;+/�]��S�x��g�O�͌ӡ��"FZ�;V����u>uT�̯B�Eu�죜�"�1<A���!���X�U4;��������h������^(���*��^A��*�d���kM*��J/hmoo��շ��^Y�]_[�ߖ��=��C��)��ȪΙ&��4?�BK;Q��Ċ���F�˰����##�<0��x�!vw4�m�d��q��j����G�k���$Ql�{����R~7��RY��P=��\���x'�gs�H�֎��5�ׄ���߂���T!�:��Φt{"��k��;P���
��� N 	%�hYԯ�p� ��
^U�,�Q�)�>�[v���[�X��i�/cV%���,����j�&鍩���sC��\m�Wz��_d�U7�s�֊��< @�Jd��xyܝg�7U�7l�PQ~��#0�	&D� ��];�:v;e��6�]��ZϜH=�����l��� �L,a4f�Be��$�)SG�h���K+׮]��v��B���0ߝ����9[��H��I�j����x�Ӡe)�/^H�}���ͺ�nT_q*��tc��W�v9e�Ub�Dp������ﹱW9��&���P��ͺEM�+Ƽ�1�ĎƑݽ]����)�gY��W��k዗/%���������r�꒿�t���277�rؗ��=�����g/�������Y)�7o]+�<�W��g-��W+巿���y)��\��P>z���G���r����Ȑ?;�1R"�/[+V5��Ρ6<,��>��K�0��	}��ʁ���.tR���z(��|�ir���X�KaS�s�7)�j+�ts��jd���{iHs��s�#��yg郎����j몳C�]s�����C��#������ct���W8Ƀ�23;V�.Ng�եY�ʋ���`h.��U�mt��}j�@���`p���\I�!#<)�(O��Q�|��c��"['��뺉��Vo�r��L?��(d57�p`������Pȝ��,��ej�F�@5�Z��&��۟�@�ȗ0��f��et��P��u$;;Pe8>t[pHX�8��f͹.��"�?��eՋ�rv�N����y�ąL[������
=�2����x~vT�y�%�X~�|�OE�=2<� ���/U�((	��
�F���C�Yy���� 0�GM|AhO��&eCæ&��x,u�Q5��<�P�6��±\�F���{�x5i�>^F�8�gB�� q�χ ���4���� Q������v�m�^�����|��?.O�?Մ�F��d:QZ�x	D��>]�������_����2�ث����N��vc�L��Wl(t�K2C��OXA�o��5(�Rf��b�1j��D�>b����a��v���vv":^��gEu����`���11�E�|E�~�z��G�L�e�0��Ұ��[�^�b�����[�ճ�4�Z��0*�K�e$�^��gYR�
��ʥ+o��A?�P���:��@~���w��%}�� ����ظ!��G�Rv�tc���W���$���F���о�5ێ���<f�����GEc�)����PғJ�E�q%3V�]�R{E��%/�����Q988��֭Y�ώ�����Fxcc�llnhl������%�͟�2	��(2G%u�,�Ҭ~'�m�U�s����RN˵����~����O>�-�pR��˱ƺÃ�a�6[�)3��Z��p7����l��I�J�x}e$>��v(5x���n����c)S�wnBGF��蘦�Q%�'�pFy)�1�G���nF6wv5��{���w�n�?i\��F�J�bz�B�ŏ�C�+�
� �%�_8�je���r�_��0����wyDn#��:�.�Fȱ�n"D+oB�N� 6N�A��cu!���XA�e�1q$�+��M$vث�_'��O�y1bD�y������4���H�bS�)C'��4�@p;QȽ���z*�m��16�ܲ��8��{����sv�}rx��Q��6�������3��[yq�*��r�l�W�a�/�����;���6y�aqqNq��Q-s�Se��*3F�o����Wc���QFXq����#�aX�b��ܤK �Lt@^<+S3Sejz���+�G�<�|Y������~����_h@�Єu������w~V<4�z �Vi���P���)��@ۜ�B�*VH��W[I�+�E?
>~�w,X��+�<�����*S?�cE���o�/�^PLeZAT��E�(�~$}a�E%?��bs?'LЊ���fI� �؈g��4]��G���C�����h[=5WT�cV�|rC���'�f
�ٞ�Chy�7�e�)��I���F>��P�kxq�������x�g�g4,�/�����:6�e���q,��f��qy�(�p�Ɨ�<�Z?�9>a�Q����	��A�Y@��(WXɽ$z5���k�'qt[X83uzn�,.��bY��P��ʼ�P�+.��׮��7���ׯ�kKKenf��\�(��J!�!B��V��x���GV[�����*٣G��>*_|~�<��f�}�ZY�x�� � �Y��HC�o���mOd����s,ZUl���<]���Zy������Vy�8>W�f�5�ϔ�8�bt|����*�{'euc[�Y��Ս��*�]4�:�vM��Rj��E�Ę�A��h*6��竕Z�H���ݞ!;P��b�� �ς�J �Ŧ��-bQfu�3Є��ڿ����h�xt�[J��3�ㄉ	�&`�16zş����4��!pT��f�%J�y�N_��pjx8z<~�L3�����Ԭ�a���$�_x��=��f$�[s�	J��2QRp0bRh�Nj�nC�^�P��� ۍ�lH���.����r��K��� �`P��|��_LҞ8���Ǡ�� �^����M {i������&���n���_jgl��/��q�+�G�Nӫ�ellH�d�zm�ܾu͟ �"k�@x+�(�3���|��uM
7o^+7nhп�I���r���rC��M���g�<hi�����Y�U[�ɱ��]�INyR��r���ݒ|�o,���)س�R-EZ+���Vb���3޹{�<��a�������=�u�ǿ��5ν\�,/_�y_0�3�5V�k�S��F}1¹��H�}3Án[�iw��}�U�6�Tl�(�l��Ȋ�1���P�eD��M��3�8j�8�CY!�t0$�WV�p�K>��wa�hlx�]D����pr�/HS�Qʭx���N���l���ʂĪ{5� ��«�n��&�\��2��bK��O��c�rj�mk(R5&1�Ly�ƅy���233�1�6u�~O��$hV7��n�8.���T�x�~�8Yq|bB7����^���r�|�5�Kk.��"C.�	�E[?��x,9�m��^\��u}�ܼu�ܺ}�c���mRbo\�����uA�5)�7ʃ�R@u�[qxً7��ޏ�y��q�͛os`�R>8k�ܺyC�d\�lR�Xl��?����^��qRJ/E~�L����Әvvz����W��ʳ����W0y2�X<����/���h<��a�)!u��O�����/�a���J��"�I71�eQ���ll��+[�����ً�����߬H�R�l9a�u����$=�J~�RF�y�S�Z�"��;��Q����6/iNa)u��K$��m	��L��zaP���A��ů>bC_��B�C�بΑ>�<��ϻ.��1�B67�&]~Q_ge���y��������H��,���8jaH���ʦ�����
j�\]Tg��0����rƷ��F���jB�̴:7�K#�|<nEq�pN����V�C@��pA������ˊ�.QL55�Q��>^���2�&��q)O�����=������Pp�� ]�b���FL��Y�swʓ_��Q9Lt� t�8����H+�L~a����K|¯b�;N�o������I	1�L(���<B���AJ�=_�T��B�����1}#�6�9��ϱ'�r��Ƥ!�6�S�%���N���Hyxo����?)�ҿ�'�S�͎j �����j����E.ްd��2Ս�h�Cx�d� �j'�����wϼ�n}m��o_��*���WVYq�$�#Ѽ/����p���������>���-��kbU�W5��hU�<.?:<��tIq��<���W��䷾~P���m��o������Uy�rC�WqlG�&�?�G�S`�5�K��u{V�t�'�ض�_�����J�LB{ĝ�Q��K���3��m����2���@�*;+�]善^U��A�+6��`�5� kL�G�P0�6qx�ȉa3dq�mn2�	��$��+�4� DnV��W�R��m�=����'E�dYbL5�Ư����c|�D�`@~�v�>�%a�5�m�Kv@��_ʀ�Y�קO����?����&=&rP��k�l��g���ʵ����/�?�����g����k���c�!G��h�i���9���ٍ4 �˅'�l)X��ӧo}n����5�lk�tƠ�J�1Q>r���X��=O��ę��KR�����7�xK����ى211�G��W�zb��tYʓ��?�@���bZ
��kK~Z5=ͪ3g�//����7o�?�������p~~X&&�������_|R����[���K'��|����/�6{<�G�%�u	��Q�4��tD����Q��e���?���z�V��rY���nꯌ��W��_>Բ~���G�1.�c���|KKR���(_��Q����rS7�s|V���<{�[mOŬ���}x������Iy�b����9�\U}�|�5������W���bm�s,c�ڞ������׻r��l��=(_��~�٧�������%t�K��K���ߺ�d�-kƘ,�ַ"^]Z�����[�+���t�� ��c�^^�l�W巿��g�om�hnD�E��\�ˢ�ė_~V���?������8��%x[ұ������ٟs��.+�|�7ۓ�X�eήC��%��a�f$��t���c�3�8���b��?�U[W��#�'���֝g���x�ݫr�5k��^�?����d�#{��It1��9*���
�tBO[�f�v(>
=t8j�"��� ?�!�<x�ů�/&�~(�t�weX���٨��c��9�鳢��߱r����n�&&��ʀ�AA	����֯�L�jЙ�����tݢ���u�=>9���2;ˊ�|<����ղ$s��)�w�y��j���&�K�';�{��6���=p�P�2��p<%8� 466�-��~������wo*�%�}���_�q�\��:v^�*�G��	;�C9�;��)�geM���ʎ&�?�`U@��^U�D)��Y@�ĵ�kd�z�A�K5� ��V�����*0�6P�Ic'}��:d�h��#�`�o���?��HmR|�
��������b��0{5���R��MҎ��N����6� y�=��P�t*��w$����g��$��U �&N��=x����"W��exx���X����,�ܙF�S��������1�jg�2�084�<4%JS#�⟒·�U��r[�-/S3���89��O~g5~0>�$N	'�83�1��Gб��x36ƾ�Q�;��w������%���[����۩$b��&���t�չK��?>,?�[�޻UnԱ��R"+�Ku�V�ڼ�5��h���S!>gʓV�.�������3N``���D
7۠�#O�x��E,^�c���Q�(i(�l�@��V��d�=�+ow|���+R�7�$5^�⫌���~�[�F���Ԙ��B�!����3��?ɘڰڷWY�GV�O���cN�9:�EcN��趃����~�5^+ϛ�����)�(��!c\C���eBF��~�0RD +��/�/�����K�|.���"�����}��%���#�҆l!_ �q��u���XN�.1��09�H7�l���X�=� *��'���y{��;��_q�<����3	IQ到+�o#�؎K�S��6�{�AM��σ����/{VP<��6]������-2�_�zB�� h)"�Ѱ-�Sثľ�x�ן����$������r䌉��
�j`���2}����J�F�;� Ϡ	:"u���O�~��K�.Q�p�u�-�Aǋ4j�;���c�H��� �_�W��b��0/5�g�Dnݼ�������������-�Չ�B��Ae�����}�d���jTef�=��n\��2�Adؓ�'~��
�y���%3������pt|��O^�~���M��}���yD%W�%�>�L?�(��n��L��74_Z�����Ȝ>2���=��#d�4��RP��$K�;8+�����7��Í=�jΗ�q�����&P�:�;T-��P-�& {�F�3^�����젠�4��*���T�p;��i�T�x�*/����:+�#ה��v�1�	R�-Lë��I�Y�Ե��/�C��+�Hn��N*��X�$ބE��t��e��Y���Ix�-�m��ɿ�$8o��d`�6�����$웍*+q]�N�7-���>fw�gZ@ᕥ@~�w��ba�8�`�϶zJ��Ը�����3��-��d��F�_^5��L�(o^yu�%���Z��ߏ��!�+���i�91ϱ1�\�#�	%�XdkJܼ���)oA��g�z+ �괔hNe�X4��E��b,:��F��NI9���x�a�����v�ܮ�i�-�Ǚ��!�;���7|E��h�!f�B��%�w^�d?)�V�Uf(~�o�����^��oV���a��5�v"y��~:���S!z7@l�4{q��V���M��g������!OcK��I��=��p\6���iu� �Z^//^���J&7����0�Ǿ^N�`e���t�G#�m^j�BZ��-�	��I�K�^@����<3Ut3�rKs������Դ�v������u T60�]��^9΅9ǎ���}*g�ەM�ǇRnO�O�Q��^�p��d������6�v�IV�Bʭ'S7�Kn��e�v\F�{����"�il|ܓp�K���V���@+d8��bư�-��E�7V���0��7y�ī��t�
>Hcۍ�GHlIx/����Ȋ�t�A�/����s�8�6��m�G���ޤ�~.�
�#���тT��w�}���G�O��㗓 ����w�/����0����RlܻY>yp�<|pSJ-{���`�wiQxu�\]���'G�̨��#8n\8K�/�����Մ��)�$s}�ΏtS��>Ay�A�w�B>�p��4��s�ٴ�Y�����XeO�岩�r��"5/�%�6���S�opd箟A��Y��Z\\*S�ӞpL��s0O��q..���(Y�>���8x�ޜ>�=2�خm��˻q�ʆߦ�0F>?&�`@C�]��9t�?�m�1T�����?:����o�:�Х��#eP�J������A�I{˾JP�ȉ;E��1/�~���@I#����r�_扰&����/JC'�2�_~�A͍����҈��S/��| BD��@��ȬӴb�4�t�����<"�TDzX�F�QF ���rS�5��M�M�e������*�d��~�ANG����?�����0Lǩ`�^$)a�\����J���e|�+�<�gU�@�g�:�E�I9Q]q���O��/5�h����$��i�M���Y����,���H�m	��7�(T ��Ê-�T�V���4�\-����S�̻~R�-��2��[�Wx^�yr@{y���Ԓy��}S
���F�OrQ�(*��eZ���:|���4��Mc�۬�յݲ��"��)���l�=�,O����<O��5Pm�d��Od��m�[�p��b�w<�D1�O��('�ꁕ}ŤOHN�.�/}agW��g�u���x��k�h<^_�Q�z�~h�[��qbD*�џ>�wh+얬�~[qQ?c��L��vyc]L��
7Zj`�1���=ˏ�,�h D� p�LQq�v]�fh��/IcUx��W<7�Ծ]�Ҽ[L�.�O���ի�e����_q籭
:�Ī�Q�
C�x�]��:<[�8pl�	�Qt�4�Α;EVn٫X['H�e�!8yc�-")���ΈgoR����f0�qҔ�X�>�75x�v"[.PfQ\���^�e��ζ��Q)ǊCc#ٕT�<4�I�&�=��4���)�%򆔮5��������A�I�c7�,|�suY�_L��_A�`5";\cp!�N���B���措��R\�Ǌ���:�$�6���n�/�i��{�/��יP&��L�0�l~�3�Ǽ?�;��x�/���-��O����ď�����n�-�Z��:�F|(��uL>s�AZ��ֶ:�_:(�^o��O�˳go��݁������\I�f��>��-���GF'wHJ�y��Cٖ�~xI���&�w>�}m�H�d㳛�|��@n>�{�A����}V޼=(�_���u��ZC�>�L���m�},#��I{K����ٴ;�Ym��w1�+
��J_ܐ[���m���l�ʘk&G��ؓ#�+�^���9[����jL+��q���2O\\ez�R��m���)�n�­�Q4 ��� 	 ���x(�<I _�:��U[��0�j��7x��0�-�+�#�L,�+���đi��@m;C�E�[�]�Pf	GK���"��ŀ>�rKu��s�b\۞�&[&��+�n�U&��\��i�=
��S��N�(�>�?W��|駸�����W�/�MLh>�h����U������х��eT���M���=�i�����M'n�w ��X�ζ��p���斔$>���[���k����@�6�Z��%�E�'��君����dP�q��i�r�%]ç�"ˮ��W�~x���9rV�x��v~�
s;�<��)7�(k(r��l�/646Jq}�V^�\S�m)tG2���)O������|B|[姹@u�8��dT��{n˘)���ڋ4Y�pש�~��Ѧ��Pﭛ6A_u�6���� p{�X3��x_=�ιcE��v�����M��|�g�4<?���D����%�J�}t*Y@�鐠�ɘ�bO
�>>Χ�'������VF��̘�z�֟i�4(��w
*�����)g!�|T{@���8t��`{���F���2qt�e͓�47��m�]�Ü;ύ#|�)d��ʁSC.������=/�<}��l��s�]2�\�`5:�LL�+ss�����ru)�}��c����FFƥ|̨`9"e�LNL��{�Wh�O�������`2�"��V´��(*��"��P��YyL�pW���βW-��.(�����s�c�&�ޖ���B�mOp�&O�9�W��fS����2d�V&a�.Yf*"A��7�5�����Z9�IH#y6$q����_�����+�W���[��F�i%u�Qs���y�}��e�ҩ�=zt���g����ǟ��w�f�P�y���#~Ԡ2�-�x�⊷"L��1��x�]���E�/��ߕǏ_x�4�O�&G��4@�s���W{�$�=N(�C=P(�j��H�� �ߨ�3��lA�X��۽�ۼHv��]��)G��a#�6�W^�#=ޠfG�q��&'��q\N���y�c��)ñn�����;:6�H^x�v_J�����ں�-M��JV�#7�jG^WYP��O������Ը�'L����f[�#�qH[���&ʕ����x�'��ʩ8�1�YQ����Ì}�l�`�u�cR��I�:)����(v!5���V�x�
�H�	e�=��M�+Ċ��N�ߌ��ݫ��㉓qLq��S4�*t�:c�̣J�u�Uʗ��M��|�-N�#�����L"�%�2�4(�܈�<N닜�En�(Q��RJ}XV�s&)��P>�Y����$��">�P�*B�+W�)s^�|����%�C)I~a�T��܎�h*�2�*a�?2�~�V�IP.�Z��C���6��֞��+��������)7n�gu�+�nk<	:�-n<d�cUv��E�:��U8�C^`a�髗o��ՕU)>���B�C�PG�[�>;>26\�-�ѣ�2��E���㣑E%m��m5���=�d��hߑ��X��~��͇|`a_
ܡƠ�+N
�wi���jv�Q�^a��V�xJ�6	�>֘���G&�s��6c�	H{!g[Y�����3vaʃ���v3zxt=eo�WP��Sܼ����?��y�g�6)èc�u�{qP��Ѧ��685"t8r�=l�Ff�D�CL�:[��oPƴ�0h��xĘ�֑s)�����������{����Y�3j7C��Q]�c�9���8�Ĝ�l���q�����	�v&�����mC{��*=�OP�x2¶Qn���L�������*���������NDs�&���g����Y������/^���W���N9��{UȰ*lt�&^
�7�'��Rr�PNGD	�����ڲ��K@�u�0�����ߊL9���V���ʚ�t���� ���\qƊK�|��6������3w�ꚾ8��D~��שV�K:�v*��V}�+��Z0������Pi�r��j�Íu�˰��ln�[�D���%�C&O2��@��3:0؂�Hy!^4d�H�&P��+�6=,��O�&Gک��<޿פq�/�)h��͛��E�嗟�_��#��ʱ1��������}7�X:�@|����z�ްgi}��|������V����Y�GN��2(�<Q@Y%��a���ĄFQ�{G�Z�~%u~����?ğ�Z�&{��E"?L�.#,�w2(ƑyR6�����{��S�=�l�8�����ØvÍq�Ń����i LD'2�U��ۀ1����'< `!?�Q�s�u�.�D��"GnG��+� �� ��xA�E�����Qn�5�*����΅������5�@IP,�a�P�,����[���^��2�\��^�~髚��S�[񆇸�^Em3�pOt���J��"����z�Ν�J�?^b�L���;�$)���:ϵ��
�R�e�u�xt�U��y�Mƣ���1&{/3
~$ZE?�{���/�GVH�+�e�g�yLN��>��䋛nlQnICm��'�r������H_|d��YqQ�}�-��)��kQ4�:�4-q�E����U�=;P�T�g9�zFcS}�ub�+` 
��{Ei��A��=�xI���}��W�#7�У䭯o��7+�tC�vL9�,�rK
��bTz��^Q��[^�������ɴd��7xjӀ�-�6e�Qf~!��(�E��n��5j��;�R�62�-�K����ac��~(�g�(^���7�����)�V�T�xv���N3�D��ى���i�aV��Ár���>+�~��!Zt���C�����vO�W�.1�;*����(ͮ(�&�
3t�S��!}��#�j|�|.�k���D��7�/�xX޽^�/Δ�	ՕrOa�^5+��O�C_p��Ԓ����@b��h�\/�j+R@:5�*#��&�.Hr4G�=}��}ۿ�����Cn4����fwu(�����K�������K)��_�����r�w���r;6v^fg�ʵ�U��>+����r)�����	) Rn����u:��R����\��6��le����Fa�����E���� r~ﺔ��؛!�K#��h�|udyy՟M\^��] �����2�]�.�M�L���ۃJ5��/䕝��L�F��_���2��"��)�̅[v�ReJ�s1P6�l��7ftZ5&�%�D�/�k�e����8ʼ�BGQ~�G<鄬آ�^*'et�}��N�/��_�?��'���(��\]��[����o���%�]z�<+�w��)_|��E�_.O��-�����o�)�Vٓ���Bhu&ǐ݃��,��m7��=Jy%�M�j�Vy��t��)��Ƀ��U�Pp�;҈	���%�\d
��_ihK�
�R���&�ё1�c2CQC�?�zΦ8��XY��'M�T��ɚ+��H�ڨo�x$6��c�n�d�̀z���Z�5ʁr�r�Ư@���E\׍�[���9�"n�c�8U�4��$K� +E�GXXu��!ݘ�9&��[OBQRb� J���"��P�(�����J�7�+k~\�1Z�z���msPj����u��X��#�3ڑhQ��T���nn���ꚱ�'
�g�2Y=-��۵K-�X�6�[~ʔ��w����qD#�ʶ�c���\�"/�e<�H3��8�D-Z�&�!V�d�\u�� D����9O<n"�[��;etTʭ�7p�d����S�[��W���Rxn�,&� .Ջ�x��7
.J��p2OT�!e�?
k(��'�?�s�Ę�d�im���Q�mLW莥䱂����w�;��t��U�
��L�r���2��=�P^����97��\�n(�Q�Vn�>I/��gw���^cϹ�d�LԮ�on�?a�����r�2�	�؂�ߤ�d�����C��bCan߉�Ɲ�v"i��h�$}E���^y�b*��bܦ��HwQ��&��6�qA]���1����*tű�qCD�p���ҿ̘��4b?+�W���T�皏�{�{,7�'V@WW���=F�Z!��5�R��)�!'��k8��a�����X����6%��E>K�^ƞ�o�.�=~Y����b���o��}�����T��(C�_�o��}��_�Q��1H��*y.��1F������� 2x+c�<�3���d�=r�5���+g�f֙:���4��3��N�Ҹ-��c�3!o4���#۽�����.3^$;�r������G&R�NICt*P��;]7R� ���|YN���:ѷ��D��	��vdK����
����3Ț�m� d��^���9J�� H& T>�T�2�_і8���n�䘚I�bqs�������?��Rp߼^��+_�|�O\��BV�&��5�NJi*h��n�����D%�>��|�Ȥx�7V�hw1��gBc��䊸�_�RH �Jy�hﬞ�r];�y����+ˎ��%>��Q^�Y�adt,V�Y���崔y�y��L��8)}����/u��[�4�^�}�}Rv�'-�x6+M����:e�S��8$/�����ڱ���,�4}��:CӪؽW����1503��^C�P�pi(����a2v٪�"�OQ^��¨�k�d�d�U�E:#�K ^���L�'+0�2�q�r��H�I�}��RЄgrKА��O)3�Yq�''�R��@�k�=*g���3�%��=�?�>G��Q��e+O�bL�H�m��,SYe�@(a�K���Z�; |U�2�
�$�TU�N���j�*�K*C����R���C�|�yӜ�����G:�¥��"�:F�T ��}ƝP�vd9唩@(d� ���wmDhr�4Y�-��a����C�#��ew������d%x�R�����}�G~�S7�G����sw(���?"$���{���7%(W*+Y��$���DN7o��D�xI�Ȳ�x�
d�)�m�!#�
��^�+>��� ��o�_������S��X(�� eH�X�fܫuIy
�/�XQ��~��jt��-t�j�V�[��~w
P��ʲӫ�w�ɶ�yo�}�*?P��b���� dnZ�L���^�N9H�n'�ɹ�=5�v��21Αo�=�"N���BV���0#�J�A�S�}��lӁ]vM�$DZ]$�~J�򋩚1�/��X���>�g�9m��,��M��d��nNO��9f�;���W(4~:�?�'A�8%�A�����؏aVl5�z2�DFB�0x�3���ΪX���� Y�(�D\��ֵ6�h�|iHA)�����6�-G3�r2�:2����_�42lS��J�lm��Q6{5w��O1Ͽ���|#M��U�4��1di1eL��۝�6����^���j���#S�@����&��	��D���M��M��ѵ�vޣ�j��\�;wn���t��a����������k�k��]�q���r�75=W�]�]�g��h�y�f[}�/��(���+
�A�v���l�0zr�4A��t~�v<��ӿŶ�C+�HC��(�}p���7(�(_����ꎔ�Q�XMIŜv�+�N+�U9����d����#M��S��+ϰ�`d>�Qh�$*���=nR5��1�Z��JN�T{�����)ӱ-!�X!�xt��&q��H�����q?6�1��`��i�RO���r�F���M�1�X��Q��m�+>���P>�O��+Jv��}nW��릃=�<���>��\�ZaP\)|(�(�<&�8z��[���؃�#R�����ki�]������P��������
���*���32�n�xrS'Z)��޳��Db��Pi���&U.�A�Bq�����C����'�i�'��囧v���r�-B�H����fȩHaw�
����F��N��h`��&f' �"�>T_�1��o�������� 47�QK8U-��)eQs��T�kP�	��Uc#�G�6��>�.���J�7>��|�X-e;�������r�r�i2�!;�yy��|�i�jd�~�'��n�7�����5��̒�n��ô������?�eﾰ��5��z�������wU;��1�#��5.Ջ��x\�
2F�1%<nH����ѡq���-��F��'H�c�I�t���A >��V���0��=��$�ql�\�����\�5w�`ʗ6�y��_,H�����'��X�]�~�Ql�yA�-E<I�r+e�3�������c� ��c�h ~��`2�:?D*�n��t��~�ˤ��K����^�*T�ѕ��gN�_X�t�$w����r��z���C��I��L:V(6
*�ha����^Y[�m�-����.�y(j�h�6���,�\�]-iy�J�5#�dz5T�J���)נ�VfIcf9HdZf[E�!�� ԛ
&�V�A0h��7~]�V�U�i|!giq�+�<	888�"�mmq��_�j)=���ӑ�n�)w��/���V�X����Y666ˡ�>�,��O;���Ym�����Yy	������i��F���M�p��7=.������~�,��i�aEԫ0��X)E���������P�VTō������(�H?WeG&��;�T����1�_����77�7���1�E�II�[9���˛�Q"YM$��
�ɹ�I����2�]ZZ,��3�9�I��=~�)b�/I�l�A�ť�r�F|�8>�1��h��>Gt܇��q���Y��bɩŐ�{���<;;�=^�t���'/}s��S^�J'�ɋd%ް&�I)�|�U�(Bw����Ϙ�r@�`����j�\��-g�-�J���(ܧǱ�C��-eHQuG;���T��);��I���B���חf��sS�Ug+��G�e����>��9a&ld /��(K&>G˞ՙ��2>6.���J�:�8����o+Aʳ�������?�+V�x�񃆶�A�r�����W.��Qv�)��pj��Ș�D g�� ��K�_��N�����e#���nX�m��L�nd�ڡ�L1��בK#��~���0i���i��݌EՏ���]#~(�9��|�m�IO����#wWD�3��!��	`��S҄O��=���z�*���j�!���#Ո��/�K� �;�tyd9��%e�� ���|Uz�o:��M8�FkNj{����)�F��\�o�p�K��,�/��r�:�K�#��S5f�'{��q�����J��a�|;M�N.���

ҬeA<tK?5d>��Jo�n��uT^��(?<��5?u�����18��;cѩ�W�ۅ2�������־���q�h���H��@��]�Vh@k��	�V�� ��4)'G�(\=�wBɢ�7�������J'���@�X�;`?Ӿ���c�9�V��Xr p����������<��=:x��F#D�&y�Q$ri�\�/����O�f'��h�0�^iz�WK�M҄����K���3�n��L���L#���G�N�6W�P
j�aehvv�ǖ�KI��W�c�A�B��P/�e���|y��ay��A�s���v�nY�}�|�G�l����/�̇���]��FÎpH,��`�~�'d\�B���	}"&�Oڭ�q�� C4-�Hns`���G�գ\n�-i�.{9�*�mW�PF[��vU�Ӭv���(�)G�C�q����oYyz�������ۏ鯴P�G~~4���*�1��ȍѭ�K������#O��������r���p(~(zlW)VDo�^,��\�M��[)�|:������ؓo�^��{�����v76���K#������>��۷�wMx�O"���<�����H7h{�lC8��2���Wg�8߸z��M��'RFK9e�O�8��O7 %@ڿ�,����on���?������_$��S���_�[\��efjZ�g�hV�Q&�ﾈ�����)����;7������y��?95��y���1(�_��*��噔��>�onF7�Kq��iw��H��9>�:4��r>5/NzE������E�l@-#�Q@7�k7�>��]���C���E��y-�[Fn�����W�7�S��MV���͛gH������>��Bj�?aΈe	3����r1n�4z܈�:�W옌��F�Cqb��?m+��o��>AU�PҠ�B�ſy����-�:_7�>����aA��F�5y{�$]�q��y?L��"4i`�����x ��t5�M�%;ulSN�O�:_&��:�BP��%�n��3�r#�L8�GmRv�N���ʹ#9����c-�K��Q��꘲�'{$�4+Yc�^�iP</z����EI�$����g�Wʓ�/��[�r?.'̑�+�?Ply������З��ʭ߳�'�Ra�*��Ј$W܉����N�84�دCȹ�C��"��(���6Ccbp��j�;~ �s��6�H��c�\e�v_�-{iْ���g������5����])E<��,[R��5"s�%)���b��T���m���7v~i��=XTGLP�D�iߙf�9z���9.X��Ӏ�&��.j¨�����I��l�V�W�u��a��@D:�jZ�c������0�&��)u<���$��{��eo�lnp�'�[�n�_��/�?{�	s����֖<��>}��h����~�&?h�͟bK%��,�d)�v�Gxʰ�����Y�>05�f��c�~>
�?ʛOB@a�,��9��?^,�K&I~�Ǎ}q�����yS_C�i�T��uP4�i�p��ڟ�+�TaY$3_V��7d�J�h��܇�g~U>��~�Q���Q�x��*�nV�X�O����+�|�������O�K!�Ynݘ+�c�eg��+���ew��i\@��,�o�|��Vy��-Źꏈ�\�(g��gCM��J�})��TWu6�R�\�64^l��ݭu�;-ץ>�w������g��+�}r�ܾ)zV���R�7W7��W�pw���қ
����Oʣ����%����ó����i�E�o�/��'.�jlY_c#��}�<|p���?+��������/>-��/����*�O%�5+�%�����'V]Q�Q�?��n��/>+�o�Rq^�Py~������%���g���,�`���Zˋ�_�%�I���=(�����E�c���=,�v�|��~u��O)�|j /Ty�Q����ߒ��`q팾}��x��%��#�P���6�l���O��Mn�(??}�I%ʯ�e(u���f)@���xA�v�����PPD�,*�PN����P��CIK��?�!�b~fl"��01B�m�PlaХ3-L���ȖBU$
7�1�:<�/Ao�~t���5#.���f��� K�A���Bƥܣ��^P<�TM��A�4��@����,�q#JCc;Y0(��6�j����(>L�n+jS��3�LLL��ёx
"'�)�ۧϝwڳ�Z����X�E �Ƽ��I<�
��9�q�%����[?y%|�/��o���NY� �++i���2��������*�@����uV�H��D�S�~����|*�R����$�s|*�Ll1)zR�s[�L4&;#����Y}u�r�L�e��133P`yɈo��
'�q/q��-+�[2�g�[ޡ���2�b	�%r`3����۠mok,!=�=�mO�q�H�L�G�l"}�����I��!o�o?��)~N�0�3	ы��qÌ�n��}�LLjVw�������p��~�->������6���7��Vnߺ�N:��7><|U�����ѝGq�~�My����#+�u��$+Fy��An�ru�m����L����Ǵ�E%M��p�<�
���̄�|���=w"`K׃'(?�ڿ'�nXC�:�vx8��$aJ��UU42�=�!��x�i . �M��0+�L�(�R���;�N�8�e��}��+~��ݛR��H�](��c�x���卲�vU���q��259\�_��x[J�5)�3n{g�W�2��ʪd;���(ދ^�]X���NfXY֠��V
�j����Sڏ>�-e�n�su��NIԍ�[�K�]y�R�<�4��5)�ܖ���|�H2+���Ѳ'e|{C��ڶ�=�T�@�\�B�>���&��]_*w��*_p��r+����[�T��"�䈏t�=�?�8;��>Q}��Ry��v�䓻�ѣ{������Vhy!�#��0�1�����'+[ꯇ�거0��O���R���n��kI�ɕcΎ�X��{}m]����?��B������yVc0�i��{�YpM�!�"�t$���߿�/���q��I_d����(�U.��͞|����Ug�Q��D8c@,()��:yg9�A���/�6q��M����N���<<^ل�B��0#�M�m�Wi���C8 ����#���@�݌���k���A|ʆ2jy��Ç����hC1W�t8�m9'&���Fk%J�&a����3R�AZ,�p�窏��r�p�=G��x�I2yk�j ��	�!��Q3�E�%�!��Z���ڬ�3��j,����ͭ����Z�������k,�/p��xJ���&-[��^S^�Lb�o$!%�I�h��z�)�����Hd+ {]9x��b>S�b��@��^�;�ۉ�k�����k����9��-����q�9����8�m�C�~a�O�RGdY�-b��������`���^OPj�.��!MVnѼȷ
	�������Z#��l���ȃQ�!�k���u}�Y�(զt�[�}�0��~I`�:���%!"g�.&�M�'�b��JQx��E��ɓ���)�lٗ���/�����Ņ9� ?��]_;,o^I�}���y��lnlx��e�m�=r���S_�bpY�`+@�ط����[:SL9H���T���(^qC��ś=����&�m���Û�q��)	|��i˫|�r���UNB�N5�P.	���]�����5���3�i� �+Z̸IM����~����<�|�v���x�m������GPmH��U�(�i\Q���Q#+ߪ[�^z�xg�i=b[®�wg�=Sy)�CF>K�Svn�[�[����ɱ�ea�JY�.3S�e���G*�c��P/͎����2*~�R���}un�L�8���&N�yR���ޘN����2=yY
�e)���(^�:c�U��L���a/$��b�.&�'�O��?&�O8�q�g]NO^��Wd� �1^&Q^y>��)�c���9-���7[�xbp�1��i���s���n"�[)p�F��4g�G��Ky/���(�Q�ſ��R�y%}I
�
�-"k{�ِ�q�7�P�%�z-Ov�n���	EO��j{�ޥ��u=XILߢ�j��o���b�FR���{����U�>�R��ާx���V1
��
����l�1vU��c�Ę�2aX�m�򊅥P~�;�v �RˇLzn�2����ī��ه� �/����R&��`<Bv�4EpR��0ĸ����$T$�dr�I��x��E ﬔ)��\�7
v���E�M��f��^�rUI[|�Ϋ�����S>t���Cͳ�eye�f�*tZ�NԾY�� �S&�=�7�g��?��:~�_�+r��+J�6X9��/�������+�\�v�=D��)����N�/����#��'�H
a~��')H�Y�co�
p{�}�^9�qK��2@�|J�9P���])�(�;R8��[�q�x� �Xa��ܘVb�}l	{3Yu�b�=/�I�����I����nn�R�%��Qxٳ�iӊ�
T�K�UM#r�R���^-��*D7V
����1�q
��B�ֱ��$>�� ���N��})R&y^�����:/���o��'6�����������k����A�|j��뼧��H��~�v��� �f�������ȉ�bK��n+�DD� �2+�=P��������L4-�߰��H�o~�1��C?�
eE��EIg�F�Fa�޸	l��g#.�O�Ѹ[�ڔL�� ���	�G�it�\Z�PVxZD��P�1��$%�pD�ڈ"��.�\R�=;9��ʧ�{*�}��Xʫ\+×����;�<��f�s�``�䎍�bƐ<�DQ)���6zI���339*�V�8!ErF����H�N(A�9)�|�}Fʨ���␿���	i�gV���V����&۱��g���/�q�W����J��)�ݨt��Ce�B�^����|KQ.W���_�+{;�emu�<y�|����|�Iq�m�O����~����2;=�������m�������%)�cV��V�˓���W�����w��w�>+��x���{/P��� ��Dߋ���� �0�t���	�Ca�]Rv��Y��iE���#M�I'Vp���=n�$��Bw����;΋�1nq�aE�y�sp��Q�e�H��j�(�M'���=�)����b��w"�������#��#.�#|}?~g���v����"kʂ>G]گ�Eq`d�oڱ��?�s0�P�B^L�)��Ίn$�L2OIv���zy�f͟��ؓ�t����1s��/oB�{ �Ё�Ŷ��HN�f��h�cJ�Wt>��]ݐ��~ھ��>Վ%w��.k��o��+�П�K��W(�({D���:[��I��ck0�*�:�WyT8�YEAaO�OY�����s��8��9���XAE!��7��G���j��Op�b�V�x���(���/�9VZ�ׇb�J0
-�Ŭ":n�
&�W�6���Sm���.H�d*0��Ɓ��l"t���!;���K�P�r��EȤ��� 1��1�)���D�`L0�@"�ɶ&a�+YZ��@D�}hR@F���)���&�l��@���Ξ��<'��y����G�� ����D'2M���8�
Ot�Z(��(�_C�A�f�3�(H���[|�����чj�a�<}�� ��Q�i�� �i�g�M@������}m����r�5}�q�c7<�K7m��Bfy��ik��]��7N�"/�ݻs�ܺ�25�2yｶϞ-�W��_~�ZJ[[��b{B��'��)�eN���.���l���_j,���լ�V>V3#E������T��ە��`�,-̔��'��Bw�\]���7,eZus�!Zm�@7��+[es=�����(��ȏ���Y*��c�ދfO��ry�j�lnlk;*�(�K�d[���$�,�U
��w�Q��U��8�ز*�'��|��כBMl��zr�-d�61�^�	?�-2��|���ٯ��|��weumU}먌��V�Ba���񖋵շ^�}�ɽ�٧��z���݇��V��_?)��������[)�/�˗+eM��c�^<�}�f�W��@i,
�_X����4C�޸�LC&g�]��es�<-��JyE��}��dŶ�(ù�뽍����5�F�RtVE�
I������r9��ZS�5|pYվt�/?���^�?�k؜.(��N�i�\	����_�F��}��5~�FBK_�qg:_�u��6��)����GB%]J�4y"�6`���û��|`a��x�%F&u��y��m0n��)N~�9n|����e ��#o�oK��c�W
��Ӳ�6C��D+�x�Z���W��n�/V�����H�;���^&��7�I%�n9-�n��o%
����T�)a�.�Q+�R�yA횣��W_9�����J�+R^�:��D�Ģ��u�V|Y�<��=��8HwG��i����V�xq�4h�/!2�-�Ǥ�م��H;�A����s�"�_�Y�d (�#�0 ����#�p.�]����'�g`?�Ǡ?�N<�k��[����eaaAJ�R����et4>}97;V=�Y���~���wʃ{�����Q��ǭ�p����t�EuPuڬ�^?� ������O8z<�K'ȥ0� �hg�x��7��C��Ǘ�l� ,n,Qr�|I3��I�������}O`��dj�!�� >�u����E��x��(7���t�왆�*D�?)n�*�j%[�1�sڀ�b+ (�g�g�nC�<Nu��Ӏ�{+x	�b�V�RR����8/A�����235)ER	���eф2����)��l����7��+p|�Nc7謠i������k|�[�,YY�����~����t�|�|���囯��R�B���z��X��?�I&]~�3&0nO�Υ��MO�(���ʯ��w���o���F
�W�x2��Z�m ~(���3�Ƕ���X�эȹ|�0�]��MaY)�^�C��k���o5_ly��=o�l���
��1,xzU��i��]�L4 :�Ѭ�%E��DYM�M�d�lPEH��]��(�8����87���g��8��_#��M��)�TR�=�fax�"�c $�sXS��벎1�ۂzh�|��^�(D�-eCy	�m��&�����u���~?R�ğ]����
��@�DA���$˙�S�nOp&��JIf��-������b���3�	/�)�Jєa=��ʺ��>�M������΁�!7_�w���֦�!@����Fh�`���b%/�����oޮ�Wo�����&7��'�p�#�!�pF	�_���w��������v�r�FO���Ӊ��%W�Y(2���df
���P�����c��#R���Ux��0P8Ȋ��F�ȋ,����l7���`l?�9V|���xQQ[lC�Rhyy�=�{R��M&�
G��B[l��=�����b��L�u+=�Z-�&(�2<�ƌ�KM7=��&3�t���
����ƯcXL.�m�w�s��`AHgĮXAei�4��T�4x�?�D��O�+���g��[��ya��>�V�ܞ/K��8''&��pa~��/Lɜqg��<�D϶�=O���&���"C$q���V��
�YZ�˛�ګ�d�S���mq���GE��	���+����rp�eƤ�O�	�o�ݤ��B��z[u�O�4[�����]��ǐ6J�jAf����	�|H&�Q����p=PY엩�ao[�qm�ș��у�C������r|| Ŏ����ܤ��p���
L��*����ι_@����R�6Ԧ��K�w�˜Vڥ��n�o��^n4�����_�C$�c�n[&P�P�y�uSmr�[n����Hy��}?�X\�)����w�ON?�ڏ�x�Ę9"Y9��R(]\�����,�v���W��ڲ��m�eqnN7��7Ǘ�"܎&���,%�w%�\�aU��r|z�	n�����?��O�/�^<�l;Vd9��ݻ�y��M��y�U廵��7>���ߛevvF|�4��շ|J{����8���~H��֓->	Dc��&~2mY��m���G�$&d�fr��Z�g��^������7�G���.a-PT��`��J}��ª_n0�e���3W�H�x̟.����X��Q#��j<�w�	}��+?�˃����^\D�qio���F� w]�l��C5�t{!EqqD�];2�څA:~� ���dV�= �`��^��viEKuJ�x�&��)�T���ɖdoyR�uL�:O{����ۜj� �Fr�遷!�or<��Of�����d�0�A1NoL#~`�����$x�V�0�.d�mP�~�_Vַ�K�U/t#���^�Y-k��ނ�jyG�'S�����|�I
7���}C��ڡ�/+%���2�B�V�ދ �LJ!���me��� Vo�6w����Xn������y9�Rz|����/P��B+��n�p>W-����i@d!�����G�{RvH{O�{T�$���c���{e{��+	{'�/���(X��:��J�������R|�GP,�H;HiW���(���>��h/�NPݘ�c��Zn�����@�F~m��R��!t��G�C�@�)%���T W�D�k�;1���Y���y�o�s�=���[�Mُ
_~��b����rvߐ�0���r�0�	��ɞi�Ҥ���ĢVE�	$�('奛�N��!�M���"���J��PD�F��$W'���A�(;J�u}�9����$Nԩ�'8��n��4M�8��c��J��\n0��C�o�,��������q�Ve�Bb'��M��O
X��N��嗟�?��/}T���Y��уr���23�
�~���/�7/�i������t&m��W+�)�,Ypj���G5V�81c�f���+�˰��q�թ��2%ey|r�W���7��N���)�{�X�c?���+�G;RNw���������G5���}�w�o7���z�Ҙ����`�@ț��uj�4&0���=�w]J��շV�ي �t%>[̋NQ�(0�G�.��+�����/!19�@1f�k<�P],���+�>��|�٣r��ݲ�����)+���%W`T��n��t���v�����8nI2q71z[�[�/����	`��|�B��U��цu�k���xթ
OX�+:��`L�-��0�`O>;�S��eN���i���m�n�dZvC"�V�}���G<�iy�����SV���.Ro܆����+˧1M #�'�ik}��s�cn��SI: ��'�䗣�خ�wpd����fy��&�q�7����+ōZ;F���%
�H��B�V��Ia�1��p~>��~b�⩨v'OΪ�g��~Y�����wO^�t����jY����zޣz�\�U�2��aC��e��jl!���ʿ��~�w�� c��;�2��b��#34u��,H�宓���Dƾ@^��
(��h��ug��JI�Jf]Fw���q�.�(~=�W��؛�� [!�w�۵�mU�&��B˗�N�5�I�}&~�HWf�.m�G 	������>$��i��;4��]6�(l
ϐ9W�.����h)~�Ё�O�Z���]�*�F�Ըp����C�݈���0��Cq�L�?��jRu�]}��Mm��P�8�i^�飇w}����Rޫ�ޖW�^��|��M_2�	��0�<������.�'4O9d�����W��d�\h�^�%/U�����$�#��.�����>�,����P�N��<��gi�X�H�JH])��ھ�}�!^�DSTюs%
p��҇�X��|l��n�n��f9#1���j�&ݖ/ud�p���X��s�ۓR5����r��Uݡ_/ӓS�,#��j_�8q����ڟ}���Rp?��{�z���M~��r�^ޮ���}�qc�\�\f�gʝ�w|\��+���&�T
��]�L
���B�2̸�#5�=�ط��zso���o�1)����.W��������~� �������r|�y��-��ص�=��4_ZS��u�H��
M_�qG2ݹ}S�������.�h�ԯ6ʛ7�#���dO�I����$�_|���$�s�ܸ���=*�����~Y\����/w���?/��+~�svn�<P?�zm��M��x铱b�{z����۷���{pOt�u3:���~��=����������Dt�IF�'f"!n�rbf�6Qm��� �7cZ<�d�c�d�j�����ک��+Ҍ��-��oi��ɟ|��TOHq���&�85�{$�h��k>�sx�G�V���&L�<�O�Y����4>�-�H�̘kdzNP�9e�<}>����!c ����5
�����&,���\�5L���b�c»����ԑ�����eS۬���%r�������К5�>v%= MΟ�&@��s��m��l�'��ёq!��/�Y���b&zo����̧���f:\��2�7��t?��T4l7���+�kVh���'��'/������L��e2	O:"_�i+r�nr��-�J��W��J3��>¨���-��◧�d��R�%1�C9+f�ϰ�"�""�&&qV���8 4��!��M��`[�_ �J-{k}������b&-)�G��+�LdJ�J��a�Acr�TF9�q��Dhm�W��e�5��w ��Ca`�Ft�hԃ�0`��]��0��Bp������� ��xB��^Ӳ+�l��JM�\w�Rd�[�l-x��n�w�Z�~mF���۷�Y��|�����-M���9Ufg4�Ѭ��Nݸ|%���,���ԏu7Z�N��th�nCN��,!�.[��8]H�n�L�j
20����C�u��uԏ�ϥ��_��#p]�N=�R��Щ~��q��Ҿ����9�UY��T��9\Ѻ�ĭԞ0����H���̌��wb��֍R�܊偧Sj7��e��B��4�GT��������S�R7�����M)m�[��|���r��])gsR�8��X�ݶ�V��ͽ{w˔�e���+¬��?���eJm���I���*��ݱ2��8��˾1{�zُ�}�ݔhf���y��Ub)�|��c����y�M��ny�1-�����Η���-�ʉ6/_n��(��u[�Ј�[�8��(�����Bڙ�+���\yp�N���>���kGl�x�j�|����j��s*�;�w^�$~*S�s� �W�/�ߒ�}�G�ti��8�?�ߘ�w�+�o���.�1DP4m�p_��Ƥh���G���5�Ÿ�l�'��񏨕��'PGp���0�������Z�9N�y�Jt�~��3������6^�7kZ��P˃�h���Ӡ���׼[���J���#~/T�.�K���g tҤ�"n�}mL���b蔅�9]@�0acָ@�Z7`q�܅����z��R�7?�Ra�������oX�����MŘ'��1�K�^�!�UAlE�/x5X~|)�q��Z޿�k����~�7�8�z������7+�~��V~D�/��*�YA�rФ��b��\?��L�����9-�HL���D�t�8;��Q��H���b��E2ތ�'q�Ω�Xp"���좜��k�b������Rf�h�MH;29'w?����֕Z�P�9"�JmZf8r��s�zk�GC������{���T�"�r�ʨ�V`��hP:���%������ⵃ��X�5��u\;������Bc������J@A��y��)�ڠ��w�V����μ2�\��7�|�IyG��'�9�� �"
/����+|RpďZx+�3��\/�����Y(`L篕6�.:�>Y_ʣNi=�w�>~��p��x&ȳ��LK�M��/.ݼ�2��^���l��6 g�U?�g�V����!S`�4!Wn�h?(��ߣ��]H��w�{=�ڂ��(���H����+w<`/++��A��N���V���Vn٫����O�k����8}Jc�1^��\�)u7n\����ݓ��y�y��"E�����D{E�=�w��v[f����~y�ë�R�"W���?������;����o�/����|i싟��w�K�E�w_����c� �\fgƽ�����z�	����틍��պRΈ<�͡�n�pp��yG�
���\>��>�_������V�9������7O�׿��pt[��_~~a����A��0���'~�޸nF�T��ݻao;�F�� �� �;����:��!��6��q�����e��k�moV�u���K<y=a��������е4>��wЏ��N�����$_K�����|�d3ǝ���(��d"��!��uI����>5�g�����z]d�	ﴷ���������Y�&$ڙm����n�\�. uI�{�D�����!q���V��)���U�R���S�NL���6΍w}��<y�|�Yߋ��G�crEc./��ּ�����������Z+9ؖʼ' ���'��?����R�R��\�.g��橒���W�� ŀ}
�k)!���	�)�Q�JSt��g�������.���MVϋ]����ī�n��_Z=o��i
��1Nf��Q`8B��{�Z+�?� ���T��6YF|
ȫ}��Y���4RՎA�|\��;���w�[pI]��⺊m�
���	�}����c���:�b���ـ����><k#��l��W#�:����R���V.fg�&�uM�R^�&��8&͕�o��޹s�ܸy�,]]r3\~��6qexLJ�h���<{��}�>�!���2�JӢa�:��
�n�/B�$��-�@X'ܑ?ο�'A��WM�`~nB�h���,]f�b���\�Q��k���4h� ���j\�ޔ«�4�퐔��	�������%.Oy|�nј d��&���|�%v>E`x�����%+���CY�X׀zV�g��?���&'8��1��@\)SJk~~�
.����ߦ�c�E2�%X��	RlGF�<�.��0�v��iE���o�K�|�-U�SSRb?�։/�|T=��|���W����Ј�@��3��|��hO�ԁ�?,%�E+�����O�x�tU��jy�fUc(G�i�b��Y����/�����oߺ*��S��})�꧜~�V��W�����>y�Ti�c��R�������Y��sKs�1x{sGy[�1h<�Q�T��T�h4�10n� �V�#�����g{� ��iO	�n�Y�z�4mS1�-v�1ØD"�팃Y�4?"镸�C	ԥ{_�N�|��
b�@�v���;J���5|*t"����28�5;y6������>
}R�L����Ԓ�R]��p7L(c8#VƮ��Q��Ã"��g�E�+L�Q5��U��+�<�*�A���=���7�<*��sov<Y�x���n)�i*���K��]�@ޕb\杨��-+��0�������7v�.��Vl�)��?�=�;��C��r&ŒOk{�1����I���;�(CJZ�������x�p�j0�vbEq�I:ވ�^\Vk�䲪�-�a�`�,g���ݺ�6��=��3�!G�j�Uj9>,NA�$�¤"��W�0�y�����"��`�r��ޯ"�@���qZwB�=����^@]�71��g�D�7rLu2�L��jK:W�m��Q�d���𤅮I��"�l=�$���8XÏ|�y1gF��ե%M�3j�S��bˊ�n؛��g���wn��3�(���*�����؄��215�xZ^�ؒb��o��QJ ���7����/x�ު����nX>��!D׍�E�k����WHw�e�W�h����w>k8$�Ķ�⩼��ZZ����f���"�����c�i3�	a��� ��wg�2OT�ge~vB7?��	^�3��&�#�W�������7��μ}o���iL�E(V�ܳ� ���8��xzp||\�:�W�k���"+�sR4�	�ɸŊ&G\�]Y����)�x�R<>v�/^�oR�X���^��>���[����͖��s)�w˵k���;�*�e��R���ퟔ��-��R෤LoK��5��k��ˊ��X����/?��"�rxS����Ȫ��ީO����çefv�����/����wNe,�׫�?|������_����7e������[w��{w�7��O�a)���9�?���-ϟ>��,�?��r�2�$�|l�Mޑx����]�l��1�6�h{��(�-��˶Z�L[!����4�?�-M��L%	~y�c�Wf�6� l~�#1�x.���*�߿'��b�_����¡̺�U�>"A.����@Wi[�U�#�0���0�O��H')Ý"9�ˤ�F&� ��P֠��Sl������{�cTPrS�G�FŢ ORv�v���v���.;һ���]y�'�|��������]����H�����L��B������=)���������g���W+eeuӇl��}��''(��PlC!SV@�:J��!��
JE����C�/���B��m	��Z�.��m�@��C���:p(�|�z��[��28
/Jn(���H��T!r��C,[��̄���Vm�x�X�������˱2*l�����@��6Y��A�e� ��]hd�FÐ�Q�G6��|��]҅�fB��4.c�$K��Osg��W&e*h��p�$OA��2���!�m�:���V���b�VVC,����?����%��g_���NO��,��GF����x�z��ۅ�)�n/_q\���+�����Yy�b��]���h<��-un��W1��2]������G�,@?|8���ى����>�~�0�/�:�k�1�����k��Q<R�Eڅ���-�.�n��3(;�LA^�JT#@�6�46I1�p��Ϥ���۷Y�d�������α��/���yV~x��{Z��7��(�8�6���X�q�l��c�@�Z�S{�y㺔�Y���)�Kd��"�S���kS����+��e������O�}_��B3�:���)�k��o�x��LՌ����k��
;<�8�e�'�ϥ�N�Y}��S��ٻw�Ğ���1�ǒ��[l���#��$ٖ��f]y[S�usxE
�r~�L7����޾�X>���Wl?yp���1R���������?���P>��P:����,7y���T���]�(Ϟ</������ʲkrl|�,^]P�s��%���n$�˶_��+��k>��Y�;ж����M����^������t�mL�hr\^f��4K�Z�0/0혃0�*4V6L{ �މӁ�����Jl�v�ۿ7���Of[[�ftҥO��������!b�jK���ׁ>���|;@�5��gںS��M�0�w��CnZL��:�z|�vcSн�H�u7��nTz<�+��G�X��xw��y�ǫ�ky�q/�����ē�<ueqik�P(��Z��������:˶�g/ޔRj���ڝ�+�n��j�f՗�^t8��s���bG6�oG��b���ⶔ[�׼T[��#1��r[!^Q��1;yc����F�@�.3h�U�\��J��J.[T���R�(���^oK�?�m)��������e5">��$�%td�p:��#s�V�7Dk1Wn�5�O���݄�^C8ڞ�����W����'�F������Y�C�c��	�y��dï��- �����T<)�������05H7_���Դ�1NO����	��x��R�_����AԬ=y����/7u�;���s)/�R^8��PmB��pF���椽̈́��[�N]��.�H� �G��`,J7�zh*6� ��
w����ӝ/��*�MY&M?f��i�հ��3 ���e�M]��R7o���4����SkS��i ��y�K���V8��z�~�¥2>1��v�w�ߔ��~V���ߕ�Z^K����� }h�%�m(��7p|�6�����U�`sR��ի�K:/E�=\<���xq�Ʈweey�|�����Wemm�O x���5ݔM�:c���*�<�{������V��'&&˔o�F��������SM"g�$8I�Him)��l/�SY�%���3�2�)��ݐ�zC
�u�S���|��>��n���>!<ʊ���ܽs���������e^e�V��lߊ�go��Ix�gs��1��O������(sI�O8G��e}mC��������~ymvn�ܺ}���l�K^�x�f�,����^�+úi�����47�^��z���@ۤs�W2#�iE���W��)9J�?�ׅ�V�YӰGo�~�+�������x�H{U��w������4ț��+w��0[��>b�N�.�T�c�Z������c[X�|U����u~eޭsh�VX�Ʈ]iv��M����Dn>��ۺ82�����;-|,+?������؂�6ApEc��~��%���lj�]�>{�1DJ�����c]Y�dO��;�(D����"�T6�=~�3�ʭOFB�5���
H����2+��e@!�M��Q�M#j��S��C ��D��+�=���f �]�%n��ޟ+y�Ӽ��Y�c����!	%F�����M'w���Ql�����IS��b�����Ů����Z����%�£2�S�l��a���O���:P��QE��/�s���ƭ! �tw�����Ñ��!��Z��)5��1Vц����F˨&�a�I�Н�;Mʇ�嫍��o<I���3���P��>��h��=��j�L�J��mM����x @�*a�Y��2��Ɗ��F�E�ևM�
�+�qp�{Є��Wtx5�f��T���N�V����i�:ͺ�idJ�H{�������iƉ�u�K�'���[��k�}sD�nn�&h���d�|������/��Lʓ����l�}�����,V��{e�'�er\���Rl���7�yA���>]n�����iy�r�����(͗VTG�~<�ȫ)�W��6Y�|����j˯��ɶ��:�=�蘽�R*y{������_�\�M�[Mk�d�5NYA��+�n̖����O�ޔ��e�z(�#٪_o�-��YQ���R�-�O?�[>����Kn�uT�p�.'�4�O�x�S��!��O�	ݔ��e~q^�q�C��䑕ﭝ-��ڍ��&G���}��
�՜'ϔ�Wo�|s�q��Q�g��JԦ��ad�Z���.�C
�6A[�.����h�A�� xbP��P�sZ=�fh�����^i��e�!�5е,������~��O\rnL��Wt>\X�kK��)��O8JͿ3	�kX�?���3͈�gN�5t�(�`�f`V{7��t6�)MG�*�g��_�#�� �B/�D����@��0��jxAD�p�v��D�P Ï��迼����/����+��Z��nh�[��.똁��_���%>��X(�(�[��ǵ�]�[+�IwC��MyԼ�b�F�\?Av���KVl%�
�r;r%�ۿ�����нrA�P��qdR�����4��c���3˨�>L0�0U�I�^�����1	�Qj����Cw����.i���)�b!��+:[��RU�� I>�ߔO�(���G2u��T��Y�]���\�`2b屿�$�J�L8>����
S�|3�7�0�_i�k�.�j6��j�|�6���x�|^V&�Lħ��.������ڢNpZ�,�'Oޖ�.Ϟ���§@9z��*�E��o�s�t9'�Z�OGц,b�W�n��Cf�0г���$�eqӍlf٩�.F�1ӏ��Ε8��|��D.�7n��+���3�zO;
D#�H?���jj�52�=�������/�Jv�O��TV�I!�-��9����}��7o6�:@�����r]��=)����yƒ���xw˫7+���O���*Μ��%٧��6����6G�<}�\�ɟ�ޟ�����
�}������om&�	������^x+��Vy7��9�~��|���巿�]��o�*������o������H�u)��bGH9��T}z�|��O�g�}Rnݺa�����Ǥ���{u�=�Kv��-���ûޣ�s����ӕ�253�r�Y�����I��/0Чg����X����*���I�̛���g?��_
�|�����J7�_+_/^���)O\�p�C��Fe�b��~�D�1�4m�6�/Ǩ�N�iG{��k��D�'�X5��5��j�q���&����4-�^������{�ï�祏��h �1F��cS�s�T�un�_�L�#^-~��u �JO|H�>D�B�a�a@&bVW$��B��C+�m�Y�!��E��#�}
�mPv�o��J�?���'���3��H��8x�.~ԏOK��\t,ŉU�p��lK�����d���lK�c(����͌�<�⋲l=�	��J"J-:i��&2u���d�^[��,�,ѸPn��Ӹ�ۿ�oK�m?�!7C8S��~io������FW+)*�C�HW��4���5�ǋCh�I_�;õ\h��f�����'}/��Js�,�4�b����ʳ'܃B��(��9�����sB������&�h�M����0e�vyF����wx��G��ǰl����)��G��8jD��9c�M�|u�u}�@
ʶ�0z�|��z�Z�V��AX�c��;��sn�\������QywY5����H�1�Xeo��ٻ��A�:��[�(�dF�ˑH��,æ\��E����l����k&����v��W�Fk����\!���&^.��2���i'(�|�����޽w�ܸuM
�t-犻�w"%���[VV�<Sߣ��R¤�޼^�޿S�������{+�������}49=�t�ݸZ����M�������D������������L�;������re��LIYT��f��^��OW���1�WFF$+�ǚ�D�Y�6�$�N��ޓ<j�g���ڍE��fy�������̩
ܼ����U�<��<VF�g��/
���7˧��+�ŋ-*v!}T�]t<MAa^XZ,�Ӛ��|���w ��ۉ21�r;a�v����LKƅ�K���U�8W�c�1����^�-�?~�Ǚ����9Y��qd��`�R�!�V��>��^@�G�?���ڡQu.�@���aoe�E����.�CK��r�x!- ���+�w��w��E�soP^}i�!�<��PţY8�/n*�fzƴG��Z� �3@�v�X���x�����@O����v��/����aԧi�������MVR�_��b7�
�t�\��e[�(�˹��47��z�n��˱���=n��(�؏���V������s�|��j��S���V͏4C�h�r�=�]���\��r�w(���kb�L͑�0�-v��kZ����{v��a$�����Bh*]�^*��.H*=`.�0=� ��U��-�#,ܘ���Ҵ�9��N���[E�	Z���Е�b�����a�Jk���7.����[yF>h"��|�+�E�AG�:.
2f"<�L 4�r�q�{Э�z;}�G94���kR�.+��嫵��E(�|���(�x�-	�`�
/r��Ʊ�/���Be"��g4M�5pG �Aa9dX����� ���&J �4�t*䶝v�]N�߇��q�[��F���eڔG�;nډL��yn�¿f�`�]׮��x)<A�>�q5T�:��	�Oe�A���N]�l���z��]�͞[��"5lel{ﴼ|}X�ߢ$n�m���5��f����~<>�8��HS$es��o��7�߫��MN�����(m�UM^�+�܄��8(O�����}�ύ�S{��Q�y��)S��R��<oL|z|u��mW��f{��o�����ˋ��JwLJ�qBJ�dg?j����x�����ɧ�T�,��Ɖ�N/_�U���)g>��[Ϭ��kaqQ��b�ygA��X�)o|����:���؈Wd9��:>:*�R������N4>5�#�܎4�����n&�C�׸��wT��O?}���{kk�+9�/K��Ro���:�@8��<�r��@X��dJ�lw��v��v����"G�D��w���"��՝?ф_ �B��~�&����ߋ���&��)ϟ��h�҇��|��m=�Z.�؀)����;�s�&�y%�]y�B��L!p�(���N�1襡<�f_p��~5�$���'�ŰrZ����sx6*C�'n�6v]!���(/0�I=���:��(�2c�5Q�D=���c17���'��Ç5^qB
/z;��o�U��s*�nm�<�ʦx�F�>�-��_�\?6ʧ�?�ܒ�,\�cw�H��M�J>�NFF	/]w�%Z��?,@SѦC�0ɸ���`�8�YH2e�V]�A�5�+�)��9�N�Ƙh��"۵'�^-�J�tcҴؕ;�G.̰]7��qEã?dͰ�Ob�D��_4�!�������/Iΐ���v�P'���:�e"���S;�s�5�g}m�lq���Q�,d:���y��s���ز���7
�C��Q���|I0�r(B��	���;�$O�5yD�ïPN؉��#��]�=�2�b�&���<vg=�n��/��H�!<h�&���P���>�8c�R?�_�Sg�#�M�i����h?����S33e��U)��R:G�*��S�7Oʋ�{e�m�z�j�X��������)��j]s^�vO�[��׺�B��x��Jwx���Rp��^���^i����)|M�髷��n>{Sv9�jDi�Ζ�y+�#���u�q�@�l*�W�;�'o-��e_�����1�9"�r�+m�1�Ј&V4���815Y���8gE��XUAv���������y"��+��;����W�QDQ�Q\Qf�|�����^��(�)�������N���&t]7*t�O���,4��?���k�;WUR���򻢴�s��%/�l��=0�1��o/�Պ�N���f���=9~��^�&�3��W�Ҡ�џ�4�w�`M�c���9�D��7�C'��U��ӑ;ؤ��i��<:��_�W��^҄�ÿ�m��w��]΃M�emx;?A70�y�B���o�<B���
sTS���q�(����yV�ц����.y�Y����ײ'M��ч�dѿ�O�1+EUȚp�<�j�'�ICej��/�B�',�ئ��ad�}��5V7��g��4��rUZ+Ҽ���П@�Ek��2s�X�ʚ0Ǎ��m	�'������oV�=�q�Y4�*B�T�W	ͷ���7@��	��dV��}��U0\V6˃i��
��:EE�Zx��IάO����*
1�e�WcO653�u	�hb*<��4�7g2YGjsЅ���F�F�rW�-�uA���~8t!�^YF	�r�K��.U�8����.5�=b��Lp���`����a�C`�D����ޝJi���/*����r�cҹ�Wm�]7!�-���3ŋ��LX��Š��y��A�j���rGʦvʦ.�90Բ���;q.@�\-KX�2Ub�Xt�D2��8���a���d�v�B�M��+�!F�R}d[#���#WՅ+�Dj�L*�j�p_�?&6�a)����L76g�k��r��{�`p���r���r����7�����7�}��W+ewgO<ޕ���ό��y���rK&- �����^���~�V<v�Ņ�ӲO��#�߹�3o9?�����
_${��u���W6ֶ��F���L�~��{�VYX�-����!'�p������|�Zvt�#�Q)�W����Q�|3�:��3�7���gҟ�|��b�uk�ܻ�y����7�=Է����rzr���F^������2<|I
�d�swQ&{�Q�C�s�[ ڜL&2Mj{��*�����Jy�Ó���#E{���s�f�~c�g��aosИN���͍]����d��}��p�t��c�3�8���w}���h����.0ۜ�DC��7~���p:�9mWH�L�>=$�Oc~��Z�wj�ِ~�=����|v��$���^� �:�G�{wO�.��?S|�+���T��X��B��S�0/�J�m(�q���7�tw�?�O����	wI�i?r:v3v�ʝ�1�M@�V}*�d�n8�?'u��7�,
%fu��� �d&P�	�HS�V�s5��|s���I�ap��y�s2qܿ�h��`�P�k�b���#E�O_�5��jXmRb,���8/W��ˌƤW���[�`rCT�ui�� ��Ei7� Ң��;[�j&p�ai�B|�
/B����ە��RN)�Pn�K�d� �!�+ڻ���"d v¸֌�Y+�G�����=��(f.�;�iZ2�8~����_��Y����7�ډ�YLqh�x�QP�D|�*ו&�HR�&7n��fE����Ƒ �jCBڒ[+���2���F���u�rKG�Unk���0���ԻC� �]@�
"w~����ް��A��'n���b�a֧݀��r�_]�i���#w��VrRrl�t���/��I�y{�_��ᦃ�}���O���Dـ�c|;|���NKI��QT����t/�l���m[ŗ�8����U�gF�ҵ�2;7��񒽃�c����Uvv���0o��Fjrr�,,Έ~�/(�؟-<1�8�͍���f�GY�����89�����ّ�'�_���})|��n�����W��+7p��s;�h(W����L�"L`���TY��T^ģ>�p�83��%=j�Sf�����u)�{���������W�����I���"��:کn�ﭲ�ƹ���-^�eyn^���O���>�UP�N���|���
2����v9�"�l�\)d��߅~��O���6T|\�29w9�)-O��F?i�ޅL��sz�'W���
�G�ǟ�@�a�V�9���E�-7�!l��UWP���	� 	�{Q���A4I5傢�r���I�)�֌�!w�A/��7J���w�W{��2�t�LG�2q6���h�ɨ6��o}T����|Y&���x.g�!�ʪXB�袱�-�j0ƛ^��o˦z؊r���Q�9V8���펦��7��ɫ�W*NG|�5V�ט����QeZ�r�.o���=��~~V����+�ӣ��`����.� �T��*���ť�8�E�3�1;��+l�9��d�p(�p;{�Z��3yi���i.�A�C��- �]宋��N%��{E0�Qjb��f����$�<�Ϧ��$�!k�UnA4X������G�ޞ������) ����~�A���'��xA�v-��8�y�|YFVU�r+�"P����E�u+]������E���:o��1��+�`�ٔI��.��]�,������G�UGxT�g ��ik�#n���SA�ym��T��y�~3)�K�`OL����=�?�wLyûq7ap[��z��E�1�B�G>�6*��%�~�z�Y�I�{�|��v��<�^/Ee�X�C���S�_|����S��څ�d����Q<�_ƣ���C��mNb�**��@{t���bkO)���U~��?�\��KaH2�	J�"H�?�K>�lDy���C�Wd�Ӷ)C��]��o��)���x)�g��^	��lR�����%��Q+�ʈ&V�l�r8�Q<�sz�Mf(�<Q���62��<a!�.0�5⟟Q/W\|��\~��?;S�P�ԋ�:����a�����gY�+��Z�'�sL�+��[ ����G�&t�m���!T���;���+�/I�|@����7(�~�X44}�� n��Ə>Lp�t�q�6����B��dQ^l�"g3Ι'�B��J���h*^�3a׫�ʳ�#]3���3^�kkb&�[a�r~�ሁOA�N\�w*�F��!�]�N�i�����+n��e��H�E��cϑ�j�;�h<�+�R~��"�ڃ�D�(�е�J���yɌ�[L�3��ɪ��Xp�V|�K�w�͓`�ۑ��Rn�ʍkRn������ۭ���j�b�n����⌓	2��ĉ�GS�$�
&��J�<t��e�s���f����}�J��$r婒u����T�:0����D��@��A�a�.>�`r13f2�tH�ҩh�AA��ʫ]���id(�MC�&d^u��g����t0]�S���� �i6�#��	�(@v�\Hy���&--��$*Y<1�^5�X����'�Υ�AaL������ǟI��Jm�ԮX)
���
���V�w�����Q�ip���7�
����Gz�t\��+�x1�כ����'�]�W���ʙ~9p AVL��o�m��[褡 �U;��CH�R~�H1�y�l\$��������{|t(%	��m�yiaxt�/1x�_
!�-i�����})U[�l�.;M����;�q����s|�[�N��ʱڪ��!�_���W�p}��[f���)�8�e�<�$B
��a�"����s
YuxY�-휸��*��4�!�G�&PV���',�������(K�KV|�weL�R�OQ��T�}�#R���A87�Cޘ��Z����V惬�S+��і�����2�,��]F���Y�=I?���|�5`Ѿ)�P7j[͓җ_��#��3���hC�����6;��E�~qvf��l�
�x�c��'���E@�h+N���8vE��h�x'/"t�a�Hqs��)
�s�wB��L@�0����tX�/�꡶fM�\��@�����մL闐�ԁ$�\�X����F�Zy�\m/Ck���v�5�]a��>�xC@��Lt�� �>l�����Y?����@J�;ŬG����q��|�ۺ��"���J��|����Yhs4^�9Qqo�4n�5���,�%���3��/3�#�ڒ����?������v9ˌGr�dA�&�j�V���8�� ̂���
�m�W@ZT�M	�9��+���:�
͝��r�Fc�5W�*;Ł�	�`��R	t�3pk�s@W�:|?�gi�٘? �|�d�qԐ�%��l*����ⅶ�F{����TF'���O�bv+�|� �%��EJf;ID磉C^1)��E.OȊ�|���<2�����	�/�F��+b��u�f�[��&s��q������U$..�Zmi��Qcf�kH:��~.3�6�,cpA�Qu�f9���#�߅�����l��l�~5q;�8��@�m*��/#	z�i���3��"���4p�W�Z'J��7�G��1<�<�i�=w*�Xnڏ)*�b��K[ܜ)��NyJ�}�Gq�S������2���,EP��:`e�7^J�F��D�P(��E"�2�~f�(�*g�j/Ғ�Jz�IF���mџ��s��o).陿��]#2"�PRhZʏК��Gt?��d�����AVvDK��)�hQf�N�i �wy�ۦ�!7T���8����Ƌ6�=�DHˀD�fǯ�~z�3�\s����W�_M��zE�~-D�
y��P�K%���KSf_���F�|�W+lB����$�q��u�NbT��Bt2ck\�nY(m�iWm����{��F�"&��I�E�m%KE�#���C� �l��D���ʷ��zZ��7@��r��E4�Y�%e�����[� {��˱�s���H[����հ�s`�s�q�1OA�� ����  �[�ꋥ�Gs�dяr�m��OÈ�S�����i���R�.L�������x��j'���!V��]݈d� �iqkF�A�����x+v�S��b�DGid�b4����'�ڬ�F�Ìpc:��re�@-��*a�a�t��^뻁�̙�ر��rh��)�|�d��Z�ua���{^�t�� <+� �?�N�B�r=bW�YI!nG*�9&f"w�b��&�����0 ���2IDƮ���ݾ��Y�"�Z� �yz��h�����l����P�d\��qj�dy%e���`�J�ʷ�'�F�pw��}Zi���>�6�}�x�g��8��n3�I\��M\̰G<��/vy�1��y�h��Jc/�"lz܁ a��������"e$ҡ<��j�-��K]��M�8) ��6���2F9M�[+���z�u���6�2���E^�#%�ey7�(Q6��H`SГ]�Q�ǘ��F���Y����c��� �ZN�?�=����oe�z!��.�T�����|W }����� �
<d�8]5{��n���<�(X:� ��d��t�����O�����kYX��Ƭ�?��/�h�!�m�7Za���� ���'��a�K@�pEG9D�
r��
kZ`_�������u�4�����4�Ai�W��f�%�yrh����rc6Q�f�pϑ�{��#}�ޘ����D��b�+�)Ĵ^�(�Ex�k|�á��=�c�4�w�w���x.��DW>���O��ica�mY�T6r�R��X������x�������z��* ��6���$��(�.�7�U@3^�@^i7!�\N2�̣�[��jƜ�D*O�,�aأR�X�pĲ�g��(ͼk �«���%�~�=��Q���0#�`��L�ҵaJ�'H�9�#^�m�f-c���C�W#���[�MDz/@P�brB������HxƩ(����<*a�%�;�i��_�?�9�����a��l�x�i��	��&�@�פm�y�����r�B���3��^�rw��?�R�:���t�e��0�U�A M�����-��f�>gUC-�T�д������|��>�n���(4�0�3�44��ML����v�g�1I�G}�hb���ځ&��Se�؆>B�I7Ӯ�M"aF~��1�fE��'�N%�݀�D~0I#yn"�.$h��d�iU�&AXk��}��6��6��٤t�fSǯ����_�jT�.t�2,�� ��EP��:��2���;�l����������W�?U:�#�vY��>H��	M�	�M�4�"��7b�n�핯�f�G 8=�]�=n�il���e�gY+�W�2�=�u16n�������a��I�MW��+Hrw�� ~QvM�(-h�0�>�����O���;�@�а���Pn/���2���������#�[�u'�ļ
�9��5DF��1��\"(�
���>%\���L5{.dR��t2
��N�8����4c]@�-�0L,��R�w�T(&¦��!`.�C���$y��l�7&_O�v����G���ip�/��h��-�!ZI�B�E�Hw��� jbo&���a�F
t��y!�K,GB�a���"�-3����k����sY�\*�h��^���5 H����mܤ
�����rq���`^�O�b\d`B�k�
g�^�Jn�ځt���5��_�rB�Q��uo.��x6R�.d� �s�)>��_ԟ��7$W�����
5�#���g��:��E�Mym�_�@��FQ�5�C�&ӯ����
�/�V�Qj�!�@fM?xDǶ)�2��9��x��<��@�F~��@�t� ��,�w�d�wM�5�-��K��XSo��e�5d�����aP���,�����`�,W[m �E����z������A�L���6���t;
�@�)�f�δ�<2ݖ�5E�rgPk�6��7��%��k�*��`���sX�/ev�~ ��3]Lf�?�{��E�t�X���>?�ե6�&,�Ө�M�0ߊ���c'$��D��� �u|H���]���r{���������� �������f�by�Ƭ�r�bb����x�`����Y�M����1��z)��@�����?� G�`b`��
�$whi$�ӓѻ�q)����6����z���B�OV���;�a`FGI�ގZ哷�3� V�7#�L;��x�Q�����y�ӫ�Q�a�uӀ�f�yg>}A������ �4>����
���_������E;�D�����o�L�騶�ͦɻ����t2-��m�m�F����-3�2�D��� T�!2�I����t	����^hh���^&V�X���,2]�{/�:��O���H��ؒZ_�!\��F�"�����`�
�h�*yʪ{� je��h~m&�/��ʼ`QcE^�9�Sg���I�r�-P��Oި_Aw{2�w��~�˞m��L�槲`�"?�.���/�p����r��{�MBXC�60M	#��f7��./�`�i�@܋�>�x@���A�v\��Y�@^�L� /�#�ț�#x������uu�̂s��1]va�����4�M�t+>}�	d���1n^il���t)����/��#,q����~]@���.(�8�_ ��������tQS�=���4��Ǎ�_9�i�oP��R��M+�%�T]u��.�.[p� �F<�db�˛nЕLC��XANL8.S�Cein�\�����OK��9,��G>����*�����7n�c���@9ʉ��,��v�'Hѐ��n�Mf�"�pEʭ�\E��4�ε�Q8��,o������hp�ãܡ��E��F�SN��T� J!�w��"���`�kfϲ	��ډ@|].u@
��o��`�ێ2kfh��j�B�dbc[���yid�bd�(��4(�셐 �e9��¯��Ƒ��Q��Q�_B?�7��,c�D�Ćv�A�I#����L�Eȼ� ���1�E��Zvv ��V��e|�0�d���z�$)ƎJ��VK�.�!�F8({�; ����e�s:�ݧ�v�M�����!O��4�G%l[��r2��0�Аed&����3h��|�ӎj������'_+K�V��>x,��3����#�A�+e��Ɠr-O ��O��}(�կ-�j���d������#���q	~������(���C�,��zk��ò[�p�@��
� ��o�O0�������B��T�W���~ ���abk w��|D=e�'�Ą�>�:AΏ��${֏i�ㇽ=��\&w#^qƨ�̸@'���py�*��Ƽ,�.T��������ߣ�z��L9�Zt��eC��V�G�ՏqC�LW�|�I.�A��F�M�;��)�f|j��n�T�@�]1=�Tφ>�1)�s;�D8�qg"?�r{�*����������ۥٚ@f<P9V#Qm� ~���N�ߠU?���/t5nK<E�0
��	Q�d喕[��EpO��J>K���nZ�Q�A|	��)�zg`��` Uv'�����!}��jv�U:�չ�Ɛ�ԐzND�c��?i��qX}"��ɬ�ie��|�vw�نÙ�S�4��{����޴=�:�5��Sn���.���#REy�q�'�� v��\β��Te���`�z���h �e���ȁ�
�x5�%�T.��8rpKFN:e����g&$���]^���5]躓5A�M-߸g ��`I�4+�ʗ��/R���-�H���?����r�]��Uv���̉'�o���	�J��+ R�j�8<���d�f��AȈ�΀��V��~��m!�+/^��F��!��l!9(�?i8��rkٜn���12!�"}8��l���ĳ湅�!n�WrǱ�ɷ���%��'�[fx5Y�8�+�(��#�����er�NUA/-Q��<��Б�����1k������A@�D�.�����mc	r�q7ޕO-�&oƀ�#J���LdV��-ڃ���C��i���Q��6����m�݅K�Cׁ~wD�@���i��F?��?��=�~���i�w��=�P~�ׂM��%�A�?��yK�*��
.'����8���Z����o�b���^݆~{���Qe���1�M�r嶣����������<*�*s�j{�ʭ Wn!��	 Ũ�|����� J'P���(�rcZ���SS$��dR5b��v؎i�b�ʫ�=�&^�� �̮��ɟ
��5�/��M���H�;�(HE+�hͤ9�e�[E�4C�*y^ �2��:I:��e�!/踜+D8W����Kt��wB���O��j'�֯�D�R�>h&�̛�*/_�
ë��Q=��oa�,=��d]��P���)���x�<;���2,����G�(��g�ˏ q�_�_p��v��-��g ��W;�I;�d�]:���zt�p���9^8fM�1��6~'� J+ꌟ�2lK?�7�bw��i�siA������^��m�q�F.�c�f��Єr�h�K~�	�-䊗@+#s�E��t��Ɵ|�q�d#�l��"O���Wa_�t9z,��p'�L�G�s��X=��6v���^��W>��;�v��jS2Tg��CrD��v1,|R[/�ˏ�}��ȓ�9 �2x���l	GVjCӢl{��w��ξ|?�Y��bk��&��hF{�>􏠉��/Ub��m'�d&�5�������k_�L�F��$l�R��,�<� �9������G+��)d\pL��7����[�>�6[�1�Avӄ�� 	Ȼ��4u�;�&@�6M��`q��WM�)�f��WnQnO��^��*������T��V��e��y�r�])D^�"�ܒfC���>.控����	´+��G��NT'�&2*i�,
�B����<T!�]�`w,L�5�=@�OCT�抬4��O��M��:*�
�Pd�NA����Ɖ):R#nSW���|k8h��Ϳ^
/tS�tr`��u�28��C��&�QD�� � ҷ� kȉ���h��tn�?:,Iˏ�TW�%����+6���/���=�b[�U�6���v���]@0�&�ÝC?u%���DBGI*���i���q[ے��5@1����?�o�4A�V�O3�� ������)2J���nO�d1��Gqb�!}>:1��W�&�|V.y�z�r[�,��,G��~�ɋ�%�P2k^k�����QY�p1&8���عt �@8��t���wxI����ԏ�~
�s��|��<�`�S���$=���C�#�� �����	���`P��|_�Z���br0(�={�+��ZvI%�F8�(O]l"?:c�����Q���'D���xF���v�@#i�W-O��0`%��~M|�攁���6�aY�|e8b��dH�Ė�j��>d��R{���U�� 2� �!���k���:	�-L��A��iA���<FT]��1��!��X�(:���2�zHӭ�e��Vi`��z��p����G�O*�L}�/I����a�s{�?����~��m	'g�J��X��*B�8F�R,��"�7&č��{�_#l?U���J-��)�'w�W��$u!�y��_$��
.����T��/,C(�P+��@�G��laR��߼2v�P���[I� ��e��A�h@��'���6�A��)�FNQ
)^��DIX�:]�@|�X�4���~r'20�@�Qn��K9���-�z� �v��7T�C�T+O��9�8m��h���ɶe!�~Q+��3���3̞�;r��gC�C��tL'#0K��&�i�>9T��/�@��*O���?\?�����~b|�4(zP���	���/M'x����Ħ >Yyv��5�U6�H���?y#q�����6ʭ�$�B�L��������$'�#vXP��^"�S�,:�be��L�i����j��[�ھ{):r���Sek������%��Х�=�&'�0i�9�����~ ~�s�&A��# �j�����ɴ����������/a������������O�4&���I����,?�Eh]h5�����vA�4"(��A�|�H~������<��� �C�t��!I?�?\F��@7m�4h����@F�-��e?�'d�&��c�h��е��F�Od0/9���D�)���{�gZ�]�R�U!�03~�(/�BK�����řr�?�����oV��.ʭ�g5�"*��(���G�e�J���Ǯ�aZq�/l���e"�L�d�1�H�kp���30�\�Ȫm��2фr�r(B�TW2��iZ��Q���`$ׅ���X��f��T\�̑��-e�����&l�V��Cd^:�=vE"�_�O�G��n`��i��ix�P�݅�.��B���@MGy�\���cwc��^� >���@G����tj=���]���aа%i�F������y�v�~1��0I;��G�,��i��ei����L����(0�w�Z����? �v�g8��P_|���o�6��'Ae�ig��l��s���z�Mެl�W�2�.�;Y��n��XP��Nz��rs+�8
�����ă��w���,�1+��	����rE:ͣc&d�L��� �A����ˌ�d�|�;�@%4�\�;n�k��u���}�ߎ�"���X�����?`Z;��D��?���Ɨ{�`*^D�9�@@�綪ܶ94�U�6Q;~B���E�aN��1Wak(h�g]l�XذS�X�N����v��)0�n���X�<h9�̹��
�6�{2~���U�۞��QU�����%Tn�o�������*����Kbܱ��(��ؖ�J��i(��?����4K��ǜ�̚��[ݭhnX�--�`�I���Y|�d�s�	��,���%l�swuwUu͙����;>�������#�9ofH;����{�C��<~�Oni��CԒ.]j�n��v�0��q �ĄƎ���W���_��~yy��g�s�������[�|�|r��r���_$8�R _jذyM�v*]0r��PU���H���U��hi_Q�K�;����Q�;�&��EA��7�\�$��&�9N��A�'_Wp_�}܂���Y���� @�����.W������ݢ�HcwU��A���c;���jw�䫅���t��.�_�@6rhdo)Z��wSv�����2��O:��r0G��~����d;sl����+�_����X*M�^`j<�=Sw���3�Z�}��n��2��R��1`�cZGdɎ]^^MЂ�~7u���������x��ћQj {��>����oh��:��՚���pe�*�C(���}3�7J��xg\�z��I�r3��Ȍ�3�egT�*V�q��ʝ(D�2��U9��3���Εj�kBQM���_#�<���u��'c��7er������^?D�q�<��Uj��e�r;j�C�*�`��USBc?7a�����v}r��I����T��dZ�Z4�u]UQ0�T�|`*X��持�1R@��{�G]��&�,������1�Z�0{+2U���ˢ�s�G*�[�iܿ��S�t��ܜSM�+%�d�l\��kl�]���1��M)��Ap� J��՝*k����+t5e�������B�:����:1)�ɭ��k��O�7���ۏ�۷,g<Zvp�Ieg�P{���L`�	n��b��$��,'��ae�� �:���#���/\K��=���xR��w`�	��&C����z�2�ɝD��'���?��q�����<���w�>��	����<���B�d��G�U=<���`�0���w��t2϶� y5^-sx��#�:.G0&��������s5�ɛbu�Vپ#@=>'m�6c2'��`�K@o��u
��h�+�5t�64�񀻪D�9���a��v�5�iMl`�pCs�YA�n�j?��b�?�����xt�`��v�bH��z�t��|�}�|< ��@�&Uu����0��o �-��up�M|�ۇ��0�䛾�Ryu��S�o�j��N�+�y��h;K���\��@$��?Ff���ȞGG־HgC5��=�o�4Ʀ�ʣ���������
U���Q����S�镺��_J��9�j�������C��W43�<��W�@�wcrR�'�p~G�}��FY����R�P4��j�uJ�e�5i�J`�u���
n[�_a�k�r�tTV*PUJ:��|�ߟ>_%��p�������k���r��~��pI�%��a?�O��J��Ip��|��X���BRO%ʲ�Ǭ�t���Z����h�RGw�ۋ��p����sO/�������m�ۻ���8��8['l���Ɔ����V2)�@g[�a%t W��JH~'RY�Gp[<xC�����>:�&Z�� ��m'�̪��kp�����a���!��6̾������56q�r�K����&Zܦ�Y�~�@�	(8�mJ]��n˘�C�	���H%�9?�F.2K��!en`��Y�o���zc�W�\ѓt�0�_P�����ڛ��Zw�0��S�� v������ۖYM�f��^4;3��x����UQ)�G�ǅj�M�Tv�}�w`�M����g�bM���$ȑ#dT�{G
`�4���*k�@l�t&�X�d��������k�u�|�d,@HT���,j�f����%s������Eߔ G�S�	���jRP�����T�W1EFڜ���"E_ S�@t���d�����ds�ڟ���/�{: �za��8����Ĕ�[i�t{!:u��ſVT���U��ݧ�}��O�c���-�i���y����k���h({�dެ���.�*{1D\8��/�^_�+}=�mDJ��,�m{/8A�u��$)��E	���T6׾^`���}�O���M��a���N`|8�E�F7�
�-��r-rʵ�냯9�]꟨���\ꛒؗ@6	lu=ao��ڡ�}0��@�$>�^�\��ޣ��I�ˢS��n�"æ:��_����(�}����n-Q�ь��i������F� Չ��(��|u������hQ�w"�w�i�=�T��}��hyx�:��).�Ç����Iޅ˺p\� q��6�T����O�wp�j���:��`�0�o_��;���n�BO8�mz��x��� mn���$�� �J<�;8R���X�=}�e�gh�ٜ�����sE��Dx�:~��}��n�ѵ9J�r`^U]lR/�./J���-����Q*˯L!�`P��@'�i��>����޹5�:����&ѩ��&���ڭ��=�3�d�(�Uʮ�Ѽ��	��Of0�!�kl�r��U�TP�H1�T����e~Q�B���d	�<UA@�H{�R�a�՞�/&pu��sQ!ȭ��9�Q�|�Br�#��V
7܂o\���Վ|>n�+�A�`�X�R���w&m��܈�}��IƓ�T#܃��':�4k�u��_-�D����.��'��'�u	{[gl��Im@쫂�����,{���\�L椡2I�v�
��G����֒������Us�l�z_3��׫%�P��}�d7����*����?�|�,�&^�F��Hԑy[��N�<pDF�O��8 �@�Jr��H��3��@�Q>�W���@���wOn�>�M� ���-ی��-4�,O'�\.(�d��T{�DK��@Ϳ!�t�����?�����ۻ��},�b3��֖�{��E!��U2R�QTvP[�-�ꡟ�I�	���jR�J ;y,���c+еӥ�/�v�e���)���8sp����}6�����|!;�F��uO���`���[��z�����	�&���fQB��Iuw�4Eu�� ����C�m��(�Z(���83��20ѷ��ռ���E:0|`�T�Nj߲�Vmɘh^���Zn��@O�Uv	mOV$6��)����3�hW����;h����z��d =k*]���m�m0e��&�4�l� T��}����~g��2w��ݐI����r�
5eC��LX��E֪��~�=���H�V��1�P����J�f�?y�{��%�_�-~Ɗ�]����@@%�/��"Cm�d��C/ʺi&��8�>�)R����yHl|��{�"�e��2'0KWFF�=���'�-A��T�]����n.Mk?>a~����Ծ����	~�/�VM@S���<vg�V�v��Sq�:�Ɉm<t	OYa��I��-+��5cqJ��T�#s�樉d�T���î,�~������r9�a�?@�  n�E��������I�H��� �O'c�یD&]�D�OgZ`z'�q��J6U4�T������+���y�>�	l[�����N�bB&r������rS�4m�c��nt~���&�`�S���A�
�?�6�a~�]��G�%�y�ƕ
n���M��G�[�h1�&����8Y��=1��U6Vʙ+v�E9R���Jb!t�ضh���w�<��	����j +��%%Y�����C��S�p�b���$nS��L����A����;�/#5R'!�%��{%�]�ݥ2N*������6*U2��P��7�cSω,.2�#Pv��S0_���u���-���EcH���M�������QA�f��@6ׂ�92�fa���msRoʊB'���@��ch�5�!~|xl8�[�NT�RxT{�S�l�����.��}�XXEC�����~rN���P>���4���K�a���2Z����'͸S�W�i�Ҿē�qá�{��3�{{��#�[��tIY
1E��J}j�W�i�bj!3�DN{��ύ�V�[����>�:0���,�^M�o�������e��f�gR��#G]{,G���6�}9�cu�`*��6l��u<HS�oO��0��)�~�w��̍h����A+؊'��5nK�C��@Y&k|��1�]�o�1��B(+�����ʳ0��d��H�E����m�b��l-f�]�g�i��y��.�R���%P���t8K��!{��b�,�tP%��t�S����V�I�2�j�����Q���.(U]|Ȣ>{�b%�K���m$��}U@~��%.>�~��9h�$�w��
l;���'��_ynR���p��O��=cԲU�� ����iFu�K�>f��2�.�^�t����P���ٿx��w:���(+g�P�U�Y!>�� ��:�8����Ǌ���r�@��Ԇ	�+���/ځ<�g���ҍ�_G�����_K�v�O6�ȵ<tu [/T�Kd�/G�c��5t֤>� ?�>�PO̟	`=ʩf1�G�ۧ�C���_�ʤ���yٵ�Ռ���%#D���bM��7�-G9��f�`���%@�ue��F_����Y�3�c��B��Yy�pza�l� ��;NP䶗yg��F~��hl�����4���Z�ɴ~�S����1�Q��+�M*��|U���D��`0s�[�
�)�&h�'E�;l����Ƕ�@��[�b ʏrh)rAyp����G�Q�Z��~"�=�7ټ"�<�''���#�:ͦP��we��Q/ԩ�T��3�R�|�2��̼NqdnO@��
�x1���B���Z�%�%:*2���I-6[����}B?O����L�L�vZ�ְ��1�&˖o��/�F�M~ ��S4�� E;�=	�ʧ�PL��\}��6����b���ɤ;�ʺ豥rւ,!����~�Y��y�����yX���C�\/3-_�@��`y�d����#k��	���'�F���"�����S�[sӥ� ]�1��>:��m@ˑ��Ox̉�_-?j<	l�)��kYK�sKp{��E��sڛ��_�����&�{��-9feC�F�i��6Z�O�}�|�
�=Ϣү'�:�����/��O$��k��Bl��Rp������37����_�k��[�n�_(@�w]b�@A�бDZ(� �� �(g
	���{3�s�I�x�Y2��kX˟S�P�@��~���^E��^F����;��X6� lM���3�̦�d [�� B��C�*�ھ�;5�my����ȿ.�$a݄�'���M�+6Os2>[P���ٙUЁHՠߋ�Vl1�<��n7=��YmU�cN���'h`�g��fA'��%tZ�Ǟ��Ou�'�.��`2��݄�㦎r��W�=��چ<�=�xVT�� dl|wٴWA��~��Þ��xR�uɤ�t{#p��|��*�l�yE����=��؋�z?"hX�۶���Y����:��U��>�$���X�תb��̧2�1��A��ئ���j�Ӝ#���#C��5��HƘF��L�Ӻ�c�'�����˫\R�YиӸ@��~r��&-�u����Ӹ��Ff����p�ݐi�e�G����6��V��yѡZ��r�?N��s��^�f��.[z|��!���ܐ�k'�OU2Ϙ�iw�!c�҉���f��S)'E�NN��)ѧ��Y�:A��A"r�L|�]!/N��F׬QP�҆�p�]XI��}j,���A����Mƶdt�Ni�F�i~x���P��`t�I�O���x�����b�W�,~����oݺ]��6��܄P��V8v<��'%�����m9`ֲ��؈��yu�;��zZ��<�`�c[MB�+�%��E��CGԨ�����|U0Kh6X��`Ó�R��`Tm]E��1��;ЮܐXoAgfES�\�%
dbWa�#�F��З�-�O��<ӎ:ד������	���0�I>z��O@���egL1�"��U�Y���њ��²�e��U�M�lV�rC�"����4�Z�q4c���^^�v2��v��8���l��W��b6��=l�m��9,�a���%�^߰��'����4��0��p�I����[z̋>�hiY�@ⶎ��s^PY'����1ߪ��74�`����J�ү ��c����+\N]���kL�h����]�����������xy��m�)sW�w�4��Wٖ9`���?�69��F�$�Sf�\h��}�p�XI��
�oӧn�,�����q��J�搒��h�b�k^J�jK�W����Cy����ǖ1��v�St�[�m��q*�ʣڶ�Tb�ܲ�IQ�.�ɐ�S�[O��b-�϶��$
��'�ɭ��7 ��2E@c7Jf�I���I����{��%�CY`汭خ6$��&0Yȡ[�V-&!4����\Q������ޛ��Z�ʌ(�70���Az"q���<���p��(�ӏ�}�ȓ�~bkZAw؁,�>���:	n���0%�RM��H�t�i��:-a��s�1�Gj��y/�Ex+��5�E>)��������ϖ���8�:����G�*�1]�ԙn�+�'n%�7=��.;M	�1 M�A��M�-���[�4O����U�A_ɷ�������c�1Ț�g�f�!O���m��{��1p�*�����
ؖ���N���A۶}OP&�o�!�4��>Q����U��3"+�SIs>�%����Ɠl�^�=�}�<�y:�Bّ���tQe���Ut��C�f9 5�/֕�bm�Zgٷ"UJm�a2#���_����@Ѹ�d����b�!�d;��xL�R�����"2ҍ���7 ��@��z��	�'u�	�-�T� ����� ��Mt�? ��>T���0\il#`j�"����t3�'k�u?9�ғ��:o�^tkE`���Ͳiԡ���A�L�X���*C�rH��s���6t�!R�:6u��xܦ�+ml�'`Jv�����1�u�q�Io��g�L}�{��j�
2_J���S��v��s)tqmR�6J�y����������On%�}����	u[�fB0������$_��w^/F.��m޼��@KDa�&�&&����|q,�m{�Xc{G�~'H�	#y�q�,tFNG@�O�O?r����~=Ę���}���u�灔������:�|yLh��:�@Y������(c�Jŗ�"�>�r8�?��1(�USې�i�9|�?�~vƊMg�X�K����4�84/Eo_x��Q�n܊�(�Ik��@��N>�Tl��}^ۋM���u��s���3��������vF	��qS.(٧����?��לޯ|�}�� U�.܎ ��v���槾@ڱfzR�ăAT��a�?
�Qhْ��s��?ת-�h7?ȩ��d�����(��yhm��'���s@�hM]v��m��'�v8���R�����dE��j:����V��u� ��%�$_���>�T��R�#��uC/mJMC9���z,�p�1<�.�k�t���2��T"U��ɂҪ6���57s
O��%)zh�r:!�I��\g�`	�L
�d��8'�CF�ZH�ۤ���l��Lok�G���a�!�c�y���)���U�dbD�e�	���)W�c�>^�(��~���ܞ��m��&�	b� ���]
��*41c��UA��ԫ���PҔ4U.�8x��i�[a�z�����^Y.]������f(��Cq�9��g$��}�jv������'�_k�|P?a(��$ǆ�o�ƪs�/Bh���M�®r�˾X��m�����*[n�=έ��C�hd�NH݌4����q����/kkY�d���>���*{��ݢ�`sCL!:C�H	j��3>����d�Ɠ@��8�5��D.`�PD�2󸘾H7��!�Ӂ�����;�����S�;t]�̞��N�ܹ,P�Q(�� S��Y@�Gs�=��*�GV���"�$�G�i��k��1R���ϕG;��X3�VY�4���gc鏺�o���2J�t�m�_ ���{)mK����5��J�AN@��E!�[�
�=�߀���X�puN~��~�e�K��ԷG�X4�x+���7!����|��urZ���
��QF���̇2�{�[z��M����2�m�m��cR���H��z�u[��I�Ű1��Кdm��}����t��������P�6n��Q걁J�"��+J��+�#M�u��k9�	��C|�'�йrǋū��S����"_M"�Ů�2�_K8�O������}�ܾs�~-A�QNbȚJNO���ED�+	<9���U���B=<����	���6�8A�߳�5�	��4�� ݓ\Δ~���
r��6��F䷦T�Rrde�9����i�*;u�;D�^ ���S�i�nD�.����ʴ̓߫WAX��R���g�N��p��歬�R�_5{�]'
������ͪI��?��< e�l�P�&�U�f Bf�"�C�,Y��򜪉�ܺ�B�Ö�$��&���TH`�ЦT?�i�����+l�\j�n��^`�j�E��݁�3I,��*t���_�v�D�������`[:����_-A�S�=�#uW����4���q�@�IH��]�[~�� ���h��7����.�qt� y�7�'��w�<	 ]��������2	}�̼3���'%R���^BF��1���ڟ#/�Z8aͩ�Ѐ�N�A����X�����`��ADYg%v��d�?Y��9$}g*��m/>1�<�#��,fV0��R�k.���2���u3h���_2�rl1�)�5-@^��]�a�)_���k+���h��#��J��^vp��l�&����e�U��Vȼ�u��Yo��ƍ�3%�1e�Ȫ�?��N[L�c���>U]Jw�����sP����ڠ�:�}�x��O]9��|�>Q�kS�cB�;��t<(���08��2�eV⸇��VRU�w3g�a�'^Hg��0_5tC���5�U�2�Y���K�����)����G�[!�s����.p�ێ�E�;�!��mI�7Tm{!�@�� {3�]��L~ؙ����-?�¯"���`o�2)ҷ�lat: ܪ����	WY�?�O�0�Y�����|&q�y��l��B�^	��_*#�5O�v��oj�E�x������0C��!�!)8���i̋>	i�A�|A�	�Ȝ�ey� �\����v� �]�����y�Ϝ��6���IC�U��ijd�Bh�G&X���E���2m���.� U����Y�,J'������	~в����e�l����fN�J�0o
ʩc���q`�y�j�Fpˆ�|KF�%XD����p�EDE�*� 	��1Er�3B�(r!w�diіX��ƀ(R����fz�"��m���h��mq�iǠe��`Q�{�݂Щ9�K�P�*3|覦9�K\lI��� �Oɀ�����[�[ =��0s[���2zL�6���3F�6�-�40�Fp�-T!Ě�]�Su�>�Y#�%��d��1�l��ıP�z�J��'λL'�+vT�*�A_W��8x����'���ͩ�n��Y�ڶQd�X�L��<�]o^�k�vm!����|����{�b�4f�]g�I�������!�%���¾�&�E.��HuƉ��b� [H�%�8P������7'�E���t����d޾����L��8�������J���b4^�|2�lr
CX2�t�3�S�c#��`@([�&�����#��+�i$���d����PeO��7�-;��ӎ�y�{�� pr�J�ԍ��}���.[6l{Z�%�
�&w��sj"����0�˪w`+�p�`4VyO2��ٯ���t��#���!c���	t�->��xM[8�]x����lk��ɰiD������0'�� c�z^e����`C_!�}����|�@feb�mXAu]�u�ȟ<�j��y�P�|�$�a�f(9��
�OU�u���f�vW>����v�����¾���šǅ9��� ����Zf3�Z��{>(6�-mJ�=��:���R�ִ�M�����;����=�&��uی�Y�bd�拜*r�r S�i���;N�(d;:-h����Ī��mP�������,�:�G���I�QxBM�-�
��Ю� �܎�5c�u�z��Զy�?"����:�d
�1������0���~��-��-#b��~I���m��o:�_�O,�P9�t�نJ���}n5N-l���r(���'/Y��4]hUUz�������uB��L6��YT�1q�-��j�]R2��~1/p���Hn��;�����%)�� �l	te�t����%UYH�թ��yҧ�7�[�G*]�7|�wm%3��z�8�5)Y�#��!Q|���辨*������)��u瞃[o~�;�&��I�L���j9�a����w�����I9�I[~���{ao��1�������d�WO:-j�P4�4�f&'��5Gr���O
	���@N�P̸���oY�}d�[�
N�}�r�v���&�|�j�V��Z�=�h���~�פ�b,��+�4.vL4�Lr%�:0����هe�����B>�a;<������H�Z��h���O)*<��I��E�n�����~���������=h]k���6 6Gt�����?@@���*:��8�_�֋���h���|G`T7]��ipB�
������h�gl����Ct���ro�\|�	
]hq>O�%������Nݟ]�lk+k�<�y2�ί��{(�����y9aO�H�*n�lBT�'��A[.d��� �>��� ��ּGd"$��r�q]]z��5>Il�͌�I��������擁�|7�=�S������y�jZ�x���`mu&�:������P��&R����f�
�B͞�\߹����]j�]i��@-ծ|�'�5NNK}�ښ�y-΅T�N�k%g|F��/1�ͧ���i�N�	j;�\�Y�E���y��J<���w�Q�\w|�|�C������p�Tp��	��O�mSb�Ą�od�SՑ1UІJl�>d�Ғ�< ::O��}��H+?�9�Ĳ�v�7��}�ӓ��~rpk��I���(��Z%;�����C�� �����A1;2��N��M=H�Y�t���j	n��ROծ��zC��{�|�y��;�,�2��@�g�c�-���^}:�n��{`��+��է��J�Vઈ�:S�r��A��G`����Jq���OUC����1�mLAe{l�J�g����-�7���}b��=��g�>$�K�N{���\��rl���j�&��A훋�l`=���m�*��ll�5�����FKF�� �=��`O�@���ꪪ\��9u}���n6�P6��-~k�vp���S0�ӷI��8:`3���dLr�	�c�Y[�tN���o��DדG�o�Koq�������	*�%� r{�������t������eԍ���un�v>�f�%S��Y��վ��'�GAl���QPu��:�S6�4����;��?4�AtEbZ����ȭ�1x��IG�����C!�˂��������N]]���JBOy/Y�,�u����>�t��;y��$���|��V�)B��ȕG�G�~��f��(��S���/�o���F#��kj�'2�ʒ0
n^��_��z��ۿ;8Re�%��v�40�cl�'UeR��{�pm�d1(g]���-=���z��T��
ܞ�M7�~�����z�I�_�/��ԧ�^�*��;bI�Gr���ɨ2snө6� a��nѭ6⎇������xr���[~����ϒ\i�b)�e�1X���On���!2];ֆd1J�V��t��U�}��3'�Y��9�Ol/].����NCo6�#����ʿ���⠠����2 �627�z�N��,�q{@o���59�8u�[%�Y�b�B5x5#�|O�α��ۖѢ���|�u@�����R�@��K�)�PnL�2Ý�������9c����9W��):����0ۚL����?��G��6��}5ϩ��S�����`�Q7�d_��z�G�:Vc���v��U�� ]ө뫜���o�	��As�%�N3<�����#�qi`l�����ȅB���i��Fe��L���y���Bna��RC$5�q3?���F_�[�A�f��[��E���|��BqK�heid�PE�P��-m�-�6�Ϟ@��Щ?�#�=E\ۼct��ڷ����M
n�H޸�u��!�D^�N-�hg{��$�i {���R=��63~�K�WH7�kW���7���Mgh�7������hZN瑛9���O�ͫ�� ���Z��<N��n��#�J��Q9z�FUc��Ο&H�2�JW�V��F7���N������u�D�8#J'���c��}����<�y�ۼ.��������kr�X�{A��9������|�r}	v����"T!2�We�ڐ
���KBO��h�a�S�Ρ��\w�צ�ل�s����t������vn����?�ӟ}���(����6p{���֓�d�Nj��I��$���D���!GH�.��e�2B������x+/���ց^��jy�����	З�L-����P�l�������̣�]h4���-CJ��P����Մ����ǣ��N{�@յ�,�G�ϔ��%��e�L�ŧ���	�qP��`��wY8XO	�hw�]Ǘ�l�9BG?*9a��`ɘ�#���ח�$i_}��wo��inc�k��+%c��c��|��ڞ����>A����6�]͑,�f�$B�m���=�a��s��>З|lO_�.�O|�ʚ��t(#�Py�`сH�;^eⷴ�*��fӹ��ǧ�𮶣kmGG.����'�6��ϺO~rÀY擃�dq���F_dU��s�[{�	�f�7�1v��VQ�W~��+���.$�ſ�c��V*O�졃[����w�w�j�M�  �k�Q��	@ bs28�N���E��1��'!m/V�,��� ��U.|��ä�o�N�:�����_�[��2>�֩��s���:B��t�K{�}Ӈ�{�s�F"�(2���'�~�_4�������\�5e�!ci��j1�?)-����>I�mux��!_��䉏�ă���)%�(���6�V�L��'��H+��o�;���5����^8���zǒ��+�C��5bb����pľ�g!� �Hw�[	痽�*��^�k	#��98��YBL�1�N�SkI?�qu�����@i��2�#ǲp*u�2�%�%��]�Ar��t媟ڎW�����iil�Z�X��������Q���I�ԃWwD���p�*`74����Ҋ���C>�i�l~瓄5��O����2��pZ �B�y�i��<$x��kW`'��@y��k~e�,�/y�IK��3��W�h� ��t�G��E��\yؼ�.`͵ޭ~��@R�<j�[_������r���%�.#7㇞��}�'�����4k��ٰ�m�|SY�����	O��l�d�Q8*S��p*��I�/���Ψ��w����A�������K�F��~�v�U�A/��n��`hE3���MPD�*?#G2��}-z	n���齀}o�Okv�����6��=Rȅ�B�Ip���:AK��b}�!zٳ��^.�<�J���Ǖ��̻��D?���ad�Be��0��b�������m�V�-o��}fv��~��~*���i9��5��@2��il7FH�iS����y�D3��|d;��}�����
�၆5i���o�"�宅f�%�]�����|s���|���v�v�>∆�㴴9_$���F��X� ��9�=	l�������W�(sH��� �c�*��!{���	jy��'�~�G��c;D��
+�E>
�3�~m���z4�Gk�օ�2����)ֵ)v���ϖ�~;��?1���ޜ�[�Z���˙{��uJ��d*��T�p:ʴ���tt|�+U;4,��Q�RO��gc�p`�?���[�C�/y��й���<��Τ7Y�+�R.���V��Q��6+ ae�0�j4Z�"��:�؜�MԹkyn��Kz�� �d{q�o-�C Bᝃ�RT	|��v]Ø��_��W�G�ݳ@�,o��c��n�x\�c��y�ϼY�K�|>
Oj�������\��艮R��ɳx6һ�T�K`l�>$��	+,)=J�V����EF0�֢��� ��v֚J�r�[��8�e 2��y�;�ڌ��=
GŪ�/x�.գ�FdD����Ig����L�3��	���7Yd0�����&�= ����dĘ(�/�^�
n5�/:�e���tJ*����`���O�=�خY'�A�l^K�<�l���{���l��k���Fo�Ϟ�l��^G>,��y� ����ɡ/�A�>��&d
-a'zi ���6�f�oRF&�=WC�֩jv�~�9�BrҚc�|�*���ô���+��H��>�k����Bih�CjZlL�b��j��+`v�Â	���?,i��0�J���G2��k�����vR���8PmC��(�V�Tꌮ	=�K�J��G��V��D��~�{��5�r=����XF����J��8�l����_ٜ\0֓^��&�����m�WF���m�oyJm�_�1x �z����q�5��% ��V��������W_���~���ݳ�:�Ǽ%8���d���V��:
Y6�&:�)#tb�tԏ�'�cV(���������3x�yA��Ǥ��'V������<W;�r����?��G�E�N+�p��`��8�ӄ�d�6����US��[�hZ�U�?�`���	TOr o��yp�^T^}�e(����c��I,_�v���� P�S~I.��5���,�
l�H���`~ϝ�T���rj���l��;F�S�9�3�����������eNv�N��[��?�;Bx�gC��h>"g&���	@s�o�W9"'��	�1%����2mX���I�����<��?Ϲ\��~�VC��~��$�)%�v�IhѰ��ʼ����s�r"�<��I�2�2�����y%ò����om����� �6������Ț�e�l��))�s���?Jۧ�Z	D��m4�k��}붆�fIЧdP��xe�ו&V���r�����
H�Я{���Q�-d�]�!?R��{9.bq�o����}�,g���+�y�=��X�A|=��8掵M4��P�y�LSz4Ұ���7�&?�v۴�1���y v�ʔ9�ɘ?���G]Lc���~���@�$�l��#�~��\�{�qI�u��T������C@�	���KrE�7���#}�'�m=U�V����6�0a�[(=��9�@����.��M-$�s$�L����/=�/���ݏ��w��-�K2�-�@�$��{O�S�	]6_U��p�3B:� �Z��}pkB3��;��g�Wxb���^(��j�ıZ����>5��1����x���/��W��$�ܥ���G��5�}}�)J~�ִ!D����OHp�d`; ��~.�y��;��,���*�c:��6þ?{�H�� �K��|d<����%c	2v��|���i=W�����~�H|��Zl�}��=�c�ʛD����&�'k��j�-���ÚR_�NB�a�c�(�������=�bOt��6Md��U6�7��w  ��IDAT3.~^�2�/:�y����d$�������Gf]�cG.��6�#�	
`e~��՟�唾dܳ�2��o7��G n�<����ޕ/��/�zN�|�΅E훧){p����;���Th�i� �S����=�m�ad���uZ��T��f0鞾AL�s]3�������y��~i��<����2�Hf����F��r�䞲oO�`R��e����[}x΀ L��Q)+�b����f��a�����s߶Ndg��j��'�E1��E#*6���K�݅�=w�2��rMdrd���V�����ɉ��:U��9��Y� ��A�^O&H6qק|�K�)nd���	(�FW)%+d�z~�~� ��-A�3�n����$��I���s_4�\�T7�F�xj��Q ��-��z����/��� �#��a�Mp{ey��
nyrKp�@磥�g#X�"�'���I%���[tZq쳭8ǯtP� W�	[�����s��-OQuY)�B�p�&J@�դc����l�������*���^�Ѓ]ړ
C�$��_���))���g	@o�%���4�8�St�X'�x�5�[:g�T;I9V�K/��iɷ��~>@�Φ̹�ا1Qv�b�����$�l�~��~�el�k�껽R��>� 
@������&���O�$���^�3������_�jr�)A�9e���cτE�ѯl�M���/���A;CZk�Z���G�3� }�ǎ�S[#;��yV{� 똃���4��$���,<*�y\�G��!M+M��5�����L�5}�5g�� ��v�.�����k�z7>ǻ�Tv�
���V�Đ���O����67͠r7�!UGx���a�����{�j�OA�8Sy���5��pW[�1x�}�"u:i�I��pw���1�������1����+Hf�*]�niV0�I�B�5/�^g����?��Z概[O�f(HS+Xs�.�gv��d�$�V��G�X�����,Ygc#�0���!��C'���j�E��B��]��?��?������I]��w��+�i�0q���)��wIGoǃ[:�78�O��vP�'�n�c{���C��{0�>\.��<u���������uƓ[.@B1�c:c���l�b���)\��Vf�28tQd�cv?�Ҁ��d���=a@4i����������� ���0:/Ǒ2h�+}N?At=싏;8�ߠt�)���cC{�z#鲳��c{a	��&8M�N�m�\g~��e �Ly�|����[��VdT՞$���,���Ӱ�c�/��j�3������ )���Y�z�I�#�KEHiW�:!��ʮ����kz��P0A�O�aL^ǚfP�ޯ3t����`���窦��vH�b_�f��_�O�_T3`͞_mC�eb��Е�#�}d�@9%ވ�_を��s�j�E@%*�O���~���=,7�����j��3�)�����>4���
�������ǳ�,��5<F���h*۰/7��T��fŎ�v�m��h���r,˩����y��	�~ fB����0�	��O������]Q������6
H_}G���B3��|r6t{���-���H�m��F;s̗6[D�Q*Z쓡�/���\�#/}��&h�7]vZ���{����Q���!o�Gl#�F9���&��p)���KLt6�TX|�e�SנH��UzH�F�m�S�U
����~$��������5$��b��'�;`�2���
z�:t�6��
l/]x�<������O��x�����o�c�;/�,�����[����,"����t8��y2���R�\�?f#���`��2}g��_�<(�2��*Rm�Q_8��
n��B�bqJ]�ј���Jr���*�Y��P~u���N�Gd�︭��P8�vi왡�M؎C��`��׺�����*A��jؕͯ�'�T�ea?e�NZ�u������~��h�N�`�����bs�<>���%P��6r(�g�S���&���A�%������q
N����. g����!����������a}��I?v�|.H���Ȫ�ǹ�'&_yOp;��e����#�=8ü�QU�c`} �*�Cx�
�[�����NQ�"�8��(dc��O3�J����
忾Yd�Av�DA�\a���X`�S���y<�Ů�>�9
��ͫR�Y%�_����d�����a"�>�	BN�����Z�b�]��ڟx�T���<�[�ǭ�1�Ə���ӵ�c�:E�rI�C���k1?��Ѷ�:�2�JJ�!@S���"�"v,�L���#�8Hd[P�,���C�>��윯u�mAz����dC���=�8H}��߬�1՘(]~��wq��3��Ld�����%vc>!��"���r��.��|�� ґ�F������sQ���K���SW�W^|f����}�[���7��3�`�%��c1��aaA9dge�7\������/X����KF?�u0�t���b��򢇧��5 y�����O��cM RO�8��i��n��WvS\ۻl��<����=�pL�Ɏ�.�
���a�(�1tG39��P:
qN �ς�����.IwHz��N��>`�n��d��n� 򲈜O�i���e��3{��t��A$����ԫ�;\mP��~v�Q0�)�j��\q�/��@2��PtO�i�>V�a�O�>�k����~��6٪swRCs�iM�&��:�T��޼U��c������1�~5QfuEH��`"��)�:ʩ��r��=Ecd�����~̦�ח�|�x�C��l�qӮ��cw؞�Ѝ�8�����\��B_;�fw��-�d��ba�4XH���ϣ��1��� ��*:xL�進��F��&F��G0d���{pRtcO�M["훉����{�1Z�X�>�S60W(o}��(�̵T_�:�<�����8�&z�{Ʈs�k�N՞�r�n���Y&O�ʻ}-�H{�]���zn-gRm����Q*d���+���w�Ü4M�	��_T��o�.)��v����ͫ����[~)��_O�r\�cr�ڢ�be�k�R��lV����yzKp� ��ŤMN���+�*��l�V�N|J���S�>���G)�ʓ���K��[?&�N��"�R�J�{|*0�R�+����˝�'A����	ܲ��4����ɾC�i�]���v#�s�% �l��H�,VUD��Ǐ�C��I�ᐾ�7:�d�8Q���6��nrh��3y5��?�d�>�K�N ���JW���� Z^t���G�۪�L�L�ܰ#��\,��	�8p��H�>��_Lu�d��S�-�u�ћG�ܴ�j���F�����[e��EҾ�{��p�^$�>����n��L�d���(}3�q����SF,���+6ľ-�N��x{�$e�O�f�3t�^��A�߰�w�1�����2�}F��h� ��1��c[�}�;"�l�y�A���S}U$�����T7-�;O�)�/4�q�1�Oqno�������Cc.
�ū�'���V�����T>�gA3�/h��rT����N�_'18_�\�����:�l�mO��MF��Sd�eS����q��iJ�]�jڑ�4�Qi�a�*��6r2�@m��>SEp�,���޼���W����[�w2��}��� ہ�l��CO��^m��|�-}
�pخ�f�xIܰv<��'z���'��à8��y}�A���ޒj?dҪ�:s;M���V�6�NF�Um�гC�I�~^�짧3���uU�IŴVT��5DuT��a'ڒ�����8+�;��:��%��Q���Q�͂�|���-�r�?�����B�A�M�YAs��9 ��Ӽ+'��	[��`�G^R ���朜'�����"�$��d�6�k<Gڭ����8�����e�1�Ӗ�UHLV�)T^`6���t�\��4��:�l�d���V�#�Sɒ����j�Y
<�7��{HȈ�� ���u�|�?�6��3���\�YF��`8"h�[ ��S�V9����G���c8ഐ�}[hJ�m$��Ǩ����A�V@=�!�e�hXm8
}]�q��)&����
�"����_�ə����)��`(һ*w[��IC�P�κNx�l���##(�K,��+���uX�'�Bf,Ȗ�ֲ�e'�p��+���i�7�@g�+-tc��z�D�|����j��~\�xn�r��rC��������ݟ�^��/�i�������x7�l -��4,L���_pp�P͵�V@�w^�*���2�� �9ȶ�J���8{�<��������c��d���8�"�J�`m���� }�������N��Џ��l�j��͗E�m���\��� U�X���`�r����	6�i
݌�n��$�g*z��1�BM[�b�L[0_��`���6�(۟.Y?��U�'�3��!`:��!mN#�eW��,j��	־� 5�U:W�|:6�+���x�:��ٟFuz�MA����[]t������oLo��Rߤ��o!�����Gڅ>��5�E7��j�=E�v����kq��=�Doy��Vc�qPY��?OteOl�\��-ȍ|@�
���?t�괞��"F�;#h�[��m{�"����u�	h���IY˵��9l=� 9PL�߅$�e\_BgZ����(��R��q@�?���<d�d'Lœ�k�[OrJu�s�����'���o�i��5<AG�s0���A8&r��}�����褦m����~Q��2?�H<?�YG���1���1��gu�����D�:�Jjh6l[=���s��;F��'��w�POk�/�;��O�#>�`���|�\k��=D�d�~��_Q臈�[Bt&��LC�>�N�霫��}�^Re;(}h�ʾ0#��r�|޹�e/>s��Ϳ�|���3�ljQh���ZH�6���7@�Sx!��
�ĖM���B$6� ;�.���آo�YJ�]���M2q�_z��F�����^�\V����飅J�7�J&ܪq]�n�8�v�����U�G�8�v��I?<��9u�iG���z��fN�V��F�S[UP66T�n��PA|��H��lxg�$P����hv�v�ތ����,F6aϏ�K�x6��$�A�i����p��@Ӟ��;�{�2�o�yGА�$h��a�3U3q�r��h���a��g�!oW7���J4ڛL��GI��j
nڝ��w�M�>h�� �������j�N������>����ݯ<� ��X�>d�T�y �j"��C��o�G�J������N��w�p�w��⟡�LF�L���q@׈l�޶�/f(��䔯Zg��������Ѥ��)����e�<��G�#����!b�o t�s͓�c�\_7��`������xB�-��A�z����Ol���R��X�ړ��Js:�t������T`z�&��DJ��U:���r�=O%<s�3%&.i� hI[��b�?��`��<)��к�z�&Ew?4��yͰ�'�봹��~�յ���{KV�>����G˥��kW.-����|�������l1j�t������~B[�rӮ���7�lZ���X����)*A.����J8l���z˔|�Rjyj+$�S\x����f?�-�΅���A�@�8���f7K���M�����)�&{�na@2�+� v �~rkh1�zB�f����H@�}�>��^��[��~T���~s��`��|d�������ۑ'`�[2�;E7?b]?e��J�f9�V�k��)���8�����������-�����AN�����Nt��_�.�����
�{� t֗�+��F[H
�9=�5/倞�}D����HQ=smk�{����*���?��^�ܒ�Ȃ'{�S��� ���0e_@�?u�^{ �����X����2H}U�E�c���5E�QŹ��)�`���tո��7��r�0��$���X�O��ك��W��K��O�.'���(D��8c#Or �����|���q�YO�z\_����Ujj��3�[���|���`#r��\�pT��_��3��4y]�~�����U�]���@�+4�2����#5�z����Y�) ���'��&�b�D OUy�����ab~�r-��I~
��	���!^�O쒟wEO���z�U,�=ҿHŧ䞷�	��|�v�.�"�}�|�	���\h�*�YŇ��=/<\��~iy鹧�s�P��#��rA_NξF�:���O��/,*f�9���'����p����ԯ������<X��<8��*d'���Z��8�[5=�Ytl�r.�!\��j��1D2
ѐ���ʔ�a��-��&
���/����I�u%	��F�6����[L��?wMT]�`u
U�6�Mݚ
���O���@��Z���$�x$x��� >���:����p����->¾�j*��� �r�B`!I����NEs@z�����Q�����c��G���<�1o���#���L�)O�2���9��'h�G��++�m�Sڙ��l����վ�~I#��5o!�!G��7mZ��ܞwp�����v�r�7�wm*�*�2B�[���77�<A9~l�>�]o-ԕd��b�JE�H9	ǅ�qi����^���n��UGHb�h=��qV �:7�N�I�v��>��S6$����?��94���'e0��g����U��%��-�?��7�'�؞4�<O��ݑY��d�4u��Q�n�Z��=����%��D���[I�X.49���0Nܕ������+*/(���+��༪٣:��ϭ&�t�+�(�M�%��H�M�R��5���g�W�OB{Up��p?�i��:�����Б2���c.YP�pU�u�-Д'�'�=� ���ۗ�?܆~E���W20@�"$�$����U ��_�N���d?9��D�t�:�����+t�q:]�G�T[\�� {��SyR{i��'��*�U�tg��A�ON��]LY�r��;��ť6���J��5!�%�<0��πή��O��uf�u��@7RQ��N�mj�M�y֡S����)�&��u����4����#4l^�P��t��xrk����I��J������?7�}$�M�GA-��ͷ�� g��qg���sB����tb ��	%���3�/����.L>mC�u�;cOl�D��홓��_K���̪d�jÞt0�����r�P��"�\�T�j��}�G�)@��i���֭�Ug;M�d e	LG�I]��so|fFH��&�v�.���1H��,�=��Ȱ_��^�h4�0wM�3u�*��Mb���I��n/�nzD�p̴=J[�����(���w�6P_�[P����yf�=��)����tE�!��S�?��:���������s� e�gI�X���x�!�=�T}��qy��R�\�/r>4	}tL�^�|�0�-����$s��Ê��'���@�-G�|���^� �q���?����n����%G	�!v��	:�AC�)���_�|e��=~ ��-O]�����On-q�-���N�LЫ���:Gl���#y�ZOO3���I8���X)�����l��yy���<��`,
f�������E5��x&�'�u�,��&hG�dk���3޿�:�w����$���В
��)��e�*k�
�dqN�ɟN�h����Y)h�<��t��"Z�
��q�?a3����`,��|��Z��~A741]$>�	�@XB�2dG�!DE�b��%-��(O(�X��L��ם �	a�=1���-@����L��J��~���M@��Sg��Y�4���
*c�5���o�]l=i����:�� �m�ԦZj�&iC��ܦ��_���k	X�)�
�ǂ����nC�	�>�˞d�س~�eL�-䐁"˪�y���)��9y�j��@8�+�U~���qEƏq4A���3I�`����:�����xG���tY����Ir�&r>��yt��Ǎ��si=m��&٣U��Pu�z]=�;e{A|��a�e�i5Z���?4�%|�9�'�m@6"�?k����g��y��?�sP�3E���|���S#<��`�"���<<�_�%K��*��� :���ڋ!�g�;���:�M]n��3�"E_��ܳ�u��A.��J��/�q��j��3��aBnڳ�V��(q������ϖ��/n%H�)��e`/�BU�On���w�N��@�Q��;PPK�I*U
l!*��"�T �"H *D�����xbK`{��ʽ�\��W�P�ۢ�@�Rep*̑�B��H���Lz��/g��Y��.�l#��%.����(&������]9���f�]�d�ȑ4�aVT9 U���'�@����2;h�-���khY���c�?�� 73��Wқ	�=���Ek?��?�����
э;���fh��q���Ey��>���g�c]���9$��C�OR���*'h;� nm���2JV��&%��jO(����(V��N���5m��ޫt`V>�Vfjw?���Q���R�^�+�f����l%޼.�׵�*�Zŗ���9��X'者)�����~(	�X>�/�Ȁ�;�-eG�߅�U�#m�Z�Z|�iy�)��C��x j�o�->��w��'d�[h�Ѵ#�K�PMsNG@-��r�>�~���3�u�1��_�)҆5�Ui9�1"�f^i�ͨ�m9�q�1^@���厯��w��v�b�0t�S�	�s��7�l��9��]W2����WYP�#�c||�^ڂ����Yu3PDf���s���>� y�p����Dp[���ҁ�ބ�KB�&����A�eZc�1\��=��t��~ko#v�+*�h8UjP�>	KW�"ʯ6:���ȧO�E����`#&��6 ��c,�[�^2�tړ�+|�a�qp{�y���
�����~���w�/(�!��Rhpgz�� ��e��v�߹�"!��砖�8��Ij~_�'�t�&dt���"y�jr�C� ����{��,8D��[����HNBT�E<O��Ƿ&�_�%=~B|_�v���7�p:��v!ѓa�;vF`[��1N�L�/=�|�R)�N9��� 3�WF��up �����w0�c|���ʎֹdFn�������S#c�,���\֓Լ}j<|���2�9�}��es���~%�|�mJNN9"�1�
�.�^ G�d�_`���O4�o�rL����:�ζ��vK��b�)'��L ^��&�1:�g������?>���n�Ϛ�}D��<���B���(�5Վ(*��q6�N�)��Q��5�R|m�
���:��"U���O�uN9�u=~M��N���3�
zNU�q�N�������'��S�o�C�NѕdV9��ПcZ�.���T����C�]�J4v3�o���u�wm�y���Ti�d;��Gx��uڶP=}�S?���g���W�~2�,+�"n����Q�"� �d�����T{�����Zk�����49�޺^�VpB�\�i��$ey���ǁ��X7վ��*K&�m ���L7��2ֵ0���/k˫AF�:t����QN}�x����q ���2^Q�z�h;���'��V�Op+b�2AMm�w�U�~C<(���G���n�Y���������߿��{pN.��mI؝X32ҁ�r$��:�|:]�(!`��c-F���\��x8Xv^m �*N;s@� A��Щ�A��O �-�D��]�y�T]�������@��<D���:�ZB�a,�� �k;C��9��	������H'���3���*]yI�#
�Ԝ� YB*;2���~E��xe p��~ٯ�h����˸����t��)�t�BHT��A������-�d���2|c��K]�9fJ��4�1o[� ��y����<����](��8��Ǚ�*���i~G�f��s��g��R��`_�<�?��� +��T�Mi�>نAC�2����h�އ�Wj���Z{
r���07x} �֜6$�2S���؀�6��0˙�m���t�n[�i1i���T�X=�����銧��"���P��r����%2OW����g@�/��G&bs�舘����dhn���m�?��4"Cc����[�:�=��r��l����F}�6��ts��:�"��7�@F���qp;�?C�� ���:�Xs�_4��B����AB+��@=��[��IAץ�Xw�3���ޯ��9@,��7)���|+_�� Hj�T,Ӷ˜ݿ���l\�H�*�%��^P2���I��b �=����\��'?�}��I��x'�-{�%�Ny艻�so<�U9t�C�H]&�p�n~�������xO��=?�嵄����[w��mb<�������0�2쨁q��_�������R!��9!V[�zQ�N@i��k�)���\H��B2@y����x����t���e�9&�FZ�s�1t�M����A���cp�6��V���AE?9�l���<|.u��3*l������H�A�:�ۡ��`6-� �o��f�)�#gF=�UF�F����f,�ѻk%��
�r���nFs�=�R?蝇0���<���p{�ٔ��n������ɸ<.��P>W� 9EX���D0l;�l4Ad�m��.�ݍ��2���E���f�x��m[�t4tf(Y{'h5�}z^��4�����b�T�Ӿ�N��s`s@�������
ny:b������w>6-~�2@���m�٤s98�o�g�<0�
I�6��ݟ�5J�R���4�v�����72��Sa*5��I�!�7�|�z9k�z/5�/iѸ~�I*5}��ZgLA���ODg��y3�>��Q^�^��b�^��/��M&�ݮ�miC�Ɩ�q������?+;{Mm�czN<��=�ko����j7�ݕ�nE��\'���.ݣ�ۿ���k ���8J���df�\�#���@�∋h%%x��z�w@�8�W1@�N��_tX�h7_xu=4)�6��@R�VTmuvB�U��[V���cڴq�/��?�]��`��8���+˅_���[w�> F5f�X �s���""%t9N���u��X��r���1�yxS �������M�-����(���Ӵ�(�D���_w�<46=FR!@�l�S[?�MJ`k������yc]�n����z&(]�����pV�e��J /I��[,�,nב�m\[�)��@���#c�|!?�ć[̍C|c��6ͩ�3&c~�L�Y�˰���\�du��$�Ox��z��F��&>D����놗��A�+��[�	�����]ϺZe�L?rczM��#0O-_�M[�V�VyrN�%r�d�S=u���aF����e��`��Բ��o�uJ��o�*O]n*�>���a:s�gut��B��p,�R`[��\6�4JJ�ӹ����2��dt������*`󓌺�pj��1%W9�om+�V�#H�X�̵��M�ȋFRϋ��.�4y�Os��z"��/�=����"�������TO-׬!��X��nZ�
l�I��ʳm�x�ZGc�>F��g�ǟ����e�2���!kW�+0����������<��}]fO�����9Jޔ��lt�F(uV4�X|M��O��$)��J�!���*��Yo溿@�o
h<��8ܸ�����*�N��N�,��
=ؕ�Њq�Q����~���	m��̏c�GܪG��&���Ɣ�^`�JG��:�k���hJ��)f��>��y��|�g���~%�
�y�c�2�ˊ��z#��7��e�,K�J�TW�RoA�tL�zcOz1�N��↑l�:�2V����C�tA7��qC7��7��q{�Ea�
���()�j��s������R�n�SL��U��M��	�G�Yن�ؐ���5�#*8��yB��4��������I�y-O���r�;t����M$Ys?f�6�������s~Z��n9�)k��]q�Ȏ^�	6+/"睺���(�����U��]�L��Ӏ�j[��P44y�&�Ue��*w�~^*o��n�;Ҷ�-��<C��9���C�o��w�(ZC����d�~#Q��G��	`8M9���:���r6t�C��Pi�;o�ԅk�H}�u�1Kr���U�6�-�������(���]���!<�:SkI��:�����]��S�-�唀΅f�=j��ƹl�~�����Fc���f�<}D�Le^P�`���LV剶���񕭆��J���P�}��bHOE�sW�0�\]n��2��U�EzN�+&���������!�ҳ境��˹������>���;[���N[�Ð4sUk6y��S��?���\�`@=Ic:�h�߷ժ��YнKl�lb�Z��������/�{ut�#�`TP{ο� :�����S-�w�S�;��W3��A��\���x�!�.#yl���r����6�=�V�9��7�0쐠��~�=7܍��nDl��>9u�E���r�݄a�����T~U��Pv�9��������%-9����]B�G6�1�|�V'���I�U�;�ObK˾-PQh�*D^�Ua���#�Y���<�4�-�`ua؂��W����q*��2�®o�X���j��AM�i��Qk��.�2ݥ˶4P��+3��,[l�[�|X��&�A[ֿ��_�2[�:�L`(���rC�m�Q`�	�l�λ{S̘)'�d ��yh��_�kR��X�<�p��#��=.E,��L�S��#&��Y�h �&e�Q)}3�D���96^E+���f���5�M
Ȧ�9�#�9������ȷu��A��U��P��%�@�c�������O�$���AU�g�S��?�2s��B'��s��fj�t��fE�aSگ�k�D{�I@ů?��V�c������żK�ʬ�2I�C�5>$�*$��%���������]���X�u��P��ɻ�τ]��_�����|ŃCP��$�&>�M.=���R�$����d�:������+(������^�_9���ʶ�m��>�4TT.��8�e���
N���j͎P� `��V&-X?�+~O�v��.��e⊷d�H��Mm�~ǖQ��80>,>��0�H������[��\lͦ��3�,�ѱ��$;W�Ӱ��̀�08�QOڛ��5�'�m�tB��c^��F5��'09��Ƞ��W����5�@�"��7P�3�g���_E)�b�3�!��W�'AR0�H��D#o��5D��|q�їEZ��9��*�;������~3�G��6<}l_���d�0�)���o����x�'�+M�ː⿔G�cK�w�`��j�8�]���ν�Cu���|C�ru���3(�Ǒ��1l-{]�������=��׀R3��i��HM��0j�ݪ�C�D�툽�<�z�Q�Bm�J�U=ucƁ�
69ܮ�?	fin����1�%��O]Y�U�znXK�'1�]&�LI���"��\&R����IUde�ņNQ�o�����R�4Mg��V�iJ���
��]�OmWpj~$��*	��a'�2���s`u�.���F�A����W�SP�؋v̀�_3��V�#�������>��럺��sY���(��v��@Sh�H��`�f���iM��A��@�-� uV?�E�4 �`�������M )�>��� �w8F$��fĘC���:�R��kt7�տ��E�O��S�vGqܭ��e�/>=���3)?���Pl���m���-w`�@t�2�������p'�X�i"� �2/����ց3Z�e��|[�u�a$�O�ȤCr�+Xx�� ��&�up������vd�&��j�'��e��� 2:��pUP�E��;��~���L�����sG��A��'P�c����R��_2�%4��c��U���}Z��)��I�n�� (��L�Mj�����~�N���bIv�D^2C�z�lf���f"�wJoRW��� t�= ���m�M o�H�_�A���:��mp�D�񕚜�%�J{05c�RQ�(��I��ND�7)u����
F�S`G�����Z�d���i��փ��qV���<u���?꠾���ah�ڪ� ��TQ0jf�W:ڋ��B�J��j=jn5}�,���բ�[;�h�T��M#�_������"1��tu@��F^~�Ħ��Nj)j��&�*!�TS�m�Gr�pF6��Iab�wpK�$8�,l�d�:,���4����l9j����e͏�'��]��B��z�6Ö�4���c��@������狝�u�
�͑z�U�E�n�c&ȇ#�-�H5&��<y���:hPҊ�k��%?�ʗ�4����JdV�;�)P�L�3O��$��|��'�&����
�/����Gb�un�yա/ף3��ƞ�T��r,�X+�� � �X�t��U:%�-�|~�撂[��䶃�kW����?��>��������@Jz���(u��!6H�����d����-��	ne��Q�)�@a,ut�@� ��ά2��@͏�r��'�Fd�L��V�pP�4y����v����_a�5�o}�Ƀ<0�*]>E�O8<���s'Ѿ�|�P
���:�D�6ğ3��y��߲Q��/���ܴ�n���_K��#���n@�����ID��I�CO��@E�m
��1��Q'��� D�����+�.]Op���d� �E�-p:%��9i�f��$d!�� �nh{l������J[n��h��PM��|ƕ*��%m5λd-�
�
�M]��w����$��{
�v��l��S��va���m`��k�<�j�?�6��~�]
�ͭ�Du.J�4� 5B[���ky��Ҧϕ
�!�&a>ɺ����FJ�1h�:mU ')�~���J�m��62!���T���i$i���BK�zo��!>&C���b[�#y��'{M��!]�>��Y��$�y�_:���AKCڝs��M�NW�	BgV� �j\!}���q.oY?3��#@����T�U|خ��fS`��Kf�=��L�x��w�|ݿCm;���@�3���c[��@+RJ[+��{��m]�ڟ������ܚ{4F�k�����x�.�<�=#��k>�v���}��.\��Zu�M#{b	��֟y�D3��c�
n�������O���,1���d-;r.]^��>8��<�7���?����
����	�0
����1B��@�͠P��?���= &�x\��~�ŉ<9����;�d1���o����,��I��tZN�<qL�M���e��9A����.�9��<iJ����]걫���ҳ��'@o琿�L?7(_�$k���A����?���RO"���1�,F�!վU���=r��&�3eH]F-7FZ �VlOp^J �����t�;�Y��US�nw�L+|��V�6X9�lA�j��7Ր�_#�t���d�`&�"�*�����@�2�l���- P4�e�/h0|s�J�V��kp�h�Oy��Aڔ�n1+i��?`��mCi�T����WYA�UAS�mA�IZ�~� 6�N���\��&IrHw�s{�*�m���Xm����Tl��8 V�a��1�����G�g��~M����K~�2���h��HW�CD�P5�\�(GaДG9ф|���)"��N���T1�1�g3=l����IFJ,#�B!�'p[S��u8��]�6M����jT.g��ʬ�c��%�!���%����z
Z���K��+�Ug�|G��P��u���=eZ�S�����q�ٿ�3��ⵂzz�X��1�~2ٺzN�G�-)�9�ƞ��Ob,��gͯ������}������������9�PB<;�s���)�|��/��R�Q���у���2��\�E}��X���+n{�P����˃{�,�.+�嵄����n��9�:S�"�iQ�qE:M l1��꿂]�TN����wykr�n^���?Z���� �)��'��u`��>Ci=e��Ѝ���&�	����[?%#t��
�=��\ 
�T�ڀ��D��	�=�'�qhy��mȦ+d1��S�R?���N�{h�|,�n=��$��'!y�!���B�M����g��F�.����͚�f�by"�.`%�����ׂ��a�3�*��m.�.o�������ٽ؇����?�4#����-:r^a�K,��+D0���lӡ��ɻ
lm����*rr}���W��X�G[��r����W2��l(#y��X\I�)�30? �=0���� 9B�͌3ȇ�:a����`�c��l_�n�g&�]]�:�|�ٷU���u���m��	�-O_�e�������Gb��y��"~�,�
�vP�t
�.�]3����2`���P���l;r3@O������~�S?_��W�v����6��5�?��Ue�Q��~򸁚L�5�t(%�!�����R���qʈT�hD
�]�*cM^�M������)tհ��j��)=�P�u6U}Kz�e�����k��م�d�-b�G�U�D�|֙^���4��f�?�/\�3��m��!�G:�g�E,@�I\� ���l��Nl���;��ƀy�($�!qZ��rb�N�Ё-i��ؚ�{dA�l��:��%�q{��UL��<������8�-�~�����w	n�]^�Z��"
ۨ���`��:�����[i��kp��8�E.y8 F@��V���8�:�U�B�1p`������V��`�3�O�v���A;�v`K M �:OH��V�?v[��Qy��|�0豃-}����Qv�jڝ�?��6�<��9�猋W�˕���wƅ�u*��H�\�Eͺ�Ϣ�d<�b?m��'�^����)�-PA=>��s&ԇSɌ*����Yt	n[?F��N���h]�e����I(?� �Y������M���.e�Gߒ6D\ɩ�!�E]������6��[n{x�ܰ��u��0���K�S�&�J?�n_ &���e��8�&O��A-
�N͸¾��y>�L8�xΒy��xZ*Sb{|k*l�uۆ|1�L��=�Щutڰ+#�g��B�w.T{��`�!`Z\�#+'�\���_��������Lj���f2��6`��	p?"�dq���۹���*��N,$|����|� �ҷIvCW!��0�a�|�Ǆ�,.�X*�`
�>f�JyJv�l�)�m��"���-�ɜ�T�����>��q'gv����������Q8lĦ�	e���r�҇j�H�G|"��<��{��F"do�,fCH�A�������[�'X�����S��+:�ǵ����BFɤ��2���}�r���-z����ע*���@�ܞ������%���?#�������܊��t��B��qh�H=���nыN�ly��i��tȣ�v&���NL.�qf=�����n9`��n�RƝ�#�4�m������ݛmr�ñ�0��� ��N|`�LcK��Ȕ���X���8�1��<$씸pb�r�1��y���5c�B����W��=�v)��5%�L@�|��:���ڸy�?�����$�u�4��A@�n�v@��_��Z�*]b�7��G���*���a��v�TS4LgN{�篠�,�}�.�=��%����Ď�Ӷޱ�@0?j��;WqR�*��^�Jկ�ߌ����GN'0�k��='y�)��(:o�a�BOTH�j�}]�l�|�5��o
Ƽ(<6O�J֧��٤��`�ɬ�6Ő��(2�P[�.O��un�y��
@��L�;��R��_��B�z�O�*�G@�c_�7Y������#0�oذ����IKvl-p�m�˄�-0w�PG4Տ�$U�:��*��uh���1�t����S쁌a��jچ���U����{\�kݼo_m�������kj;���5^d����FB��@q���#;E�s����;�:���t��q-klT�V�>֗��E�Jn����4�.��y@t�z@��g�Eo�~X�b�̃�Z�����el)]���]@�"�X5�}��'���Z}�}Bdt
4�狗���C��񅲧�s������d��r �P2�hp뀕2��ٯ(����y�r`���#9������c?��G�yb+Y��+�I9�(���L��1�y�I�7~��A6x�x��O+�F$�c�@�������n�(�/�;!�6��c0�+Y�U�W���K '+�2��ǐ�6�	�Z>�hM<%j�`B�Z~S9���x�/�����&��<.�hV��;ʚI$����AN#s�T|�<�*� �5/��aW�l[��t��<�/�t��������x�����Y_���������5D!�q���`k��t}Z]�z����;x/"�,�E3���˂�[v��\c.i)Wjh��m[lp<�m�ܰ�C���ᴍ3؊d���L�s�b���M�b��OՒ���m�H��Ge҃�g�^�#���+s�_�a���9P�"P"���L��6�mj��>��-��vg
Z��SK��9��q��_��M�<1���Ĭ:M"�7*���[pm����<�͐С>N��F����*�\(]]�<8ys*p��]`���൘	�#�E�wx|-g�9M�?6�]��7�2홯���w+��7͖޾>���<\��$����j�u��_�ת��؛>'�u�Bz1}�ObM�i��S���y�֯��U� A(�~��>-r�F~�s���k�Z�ѕ�V��B��!<TQK���Vh�Ȱ�������G��n��ۧ�����u�P�4 )e5��@&�4Hlw"��y�Ito'D��J�8�3xt�	��~�_s ���6�DVRg� ��Z�/�BO�82}��Ai�f��O��ɲAEz�4(�SKGC�}��@U��������N��EFH�yÆw*@2��V첏!׃1���=R:f��p�i���0�3�B����	Z��@�S�wv�k�(�8z\7=5G��O��!.������3�\5�2�/�<�����KF��Q�ˤ�iC�B9��a��g�Ǳ���&k��A�vO������vF��׾Q$�l��	)O�7��i�з�5�\������W�b�m[�;�������|h��'�oE���b���]���e��8�M8u R A֊�oʜ`�pS��W���h���_R��ՠ�n �syC�Sp_�P�I��m�����zS=G2+(�)cz�Oc|.����5�/0ϢGu��prM�>�w޲���x-��v�0�Y��b[�/#���.��X��NV5��X�}��i[�SA��Mu:��'���=��ȃ��/9O���>�?�r����)�أ��W;�O�On']��^4���:���O3u������B�8=&*��顛�J>|��7��"�1!c^͑|��(q_�}�@��-[���U���ӗ��/�	=<˿߽~e��k��9�M�#Ku;O��wp[�qn��H�1�P�T=hX��r6qp�����l�ͼ�i1���"k�����$.&W }׃R]|�K��a�;=��/_������%�X�һ1�o��]{Dol������/�8�:D�IRrG�+C�-�&�hw��cH[��c���ƒ92�* &���$�RϹ�j;H��;Gi�)sH�
��8>=@��������cJ@�yZE��ﾖ|Y�3s. y��:�<)G���l�����QC|�(%}�om�D�}�a�'��`Tk��9@�6�b�~/��YU���
љ�����3��~��Ra���L�c��-�4A�]��_����e��ů�������3�Scɚ*���Da�L`J���X���B[ȁ�B�L��4�+2F�3BG�nS�5UcCM���F�����~Nm����n
&c�5/�#-ԉs�<i#5��ι��|�����aj�i�Q��l�,��M�4x����?d�/G�ܖ:�zm�^�;��|��))FT���$��f��>@3c�i���;qD��	�J+Xn�?m���tE�%%�����4��|���X��?�o��L��0|ؖ�=6��j�1J�.��Cs�ء*W���*��%���9&�T3R�HYu�y؇sX)Veȅ��]�>��Bx尩�R�<a����g���T��'d��Uc�5u�Q�ܪ���8����������"����-�JI,����6HHZ��W�Rl��2���z��q���͗���[��Ԗ�<�h(�dc�4��*�J��f]H��ݨ�s��O��@�������ԭ���apQ�Ύ�]7k��i�c�٧�������(�?�H&	���i"_�v�F�G\���:���힌}�����GЍ(?+���*�����WHO��YPk�m��"��2�s�E��G􅖧�Ba*��P4�p��o_$���/=����Y����p��hҲ�Ck��J��,���ݧ����P�]�<�Z���E���C�hA��7O�y�,</�p��r���E�Fyd��j<�'=�<+]��@������,y�������ΐ��u�ږ�|��1O��#��o)=�c�D��Ë>�Y��.�!��1w{˅��ԭU޷�B.(�J����t�-ri�_�2��`�3Gѱb� pv~l^�� Z	|����^�=�{<P[�M��v�.�>�1��.��.�dw�[�3��N)'�J��.��s�1�E"]���6�������Mǉ�AV������
|�T���:�y�T�^�d�!}Cy���:4��pR;�s��ָrj��0�XxUq"�:��ڎa���sRȚ���3�
	h����\�^#��NZ&�V
"�4�'��uPg�]�@��,�%�I䥌���Jj3��x���]@����g>�\g�pakP�C��낯k7��3�����z�!�s���y�~n�\���7y���E��uI�S�CW�\\��ym��������wΖ�ll�,�� g�6�_2�?bL��zE�yꡈ�����&�����O2�h�U�	��t�M�R����d�/Ȼ���m�/@伐�,�Gp[w{�v��>�ah�,��@��r��:VIM/�/��q�Sti�0�N=q��~6!��m���cG��lҶz����n�!��2��>;7��
�u
g��*�_�߂L�r�/7i.{�YkCy�J�Ţ3����(��:�G�j�2k�� (��%�#0^��y{.fz�u�X7Y�d,�l>xpO���!��wU_��H-LA����-��/${�~4�*|�EuS�E|�M�s��+����`T�_��,�/�[�\=/�7����V�	��8�om�^|�\��h�z��r������K�%{ŗ��l�V��z�/Ja-`���ɐz#*��S͜�c��Gl�.�N_��&a���O���ȧ6�3���Z�<|A.�8�T&��^|L�{D\z0����~D6`�x��0V�[��Ի=s���aj��-��i�Y���7 �6���Km���D�Fx�[}�4d��w:}㣮�f���P�2��N��AWvf�s�0�'O��˖�*���f3����G�~�A6�?�^�����.���P��Ϗ7��^NKZ�y�Yiʜ�ˏ��ڣ��T�a�j\y�Wפ���Z˼�/B{|%c����3�����'����x��]d-��	B ��T��x��7�T�Z���&l��`ո(Y�9�< uEWxPq�u�˫���/�ӡ�B�Gn��ߌ�0���k�z���j�i��f�s3�C������\��sa����y;eĘ�_���%�+�9���#�}P}�o=Q��_mξQ�v���R����I�"�uա��s~����k#�*QW*Y�@���q��S�t���ECE*������+�/.7�>��M����oݺ���$���C���R���d���E�c�X:/�>�� �8�W��]�h�āYF��ǹ�c^���P�A[Sd�o�!�'��,�M�O'�F�>���������:3��/=�l_��Qڱ��U�C�n���>w��-��>�>ʒ�܏�pZBp����*uQMޔ9�D��t݌@�o0�UHIm+����JB�i�}����"�Cʙ�*hڝ	���u�ܸqey�����?�<����SO��\�^�vE&�
s^��?��r��r]�ݍ�W��7�)P���BW�<kc���Y�ͧ��"�˒�:�_�� Ķa�l�-5:����W_{�v�������
��hRI&��p�}dۯ]��<������Z^z����W^P�9���l����r�Յ�a�?]��qmyᅛ�+�<���ڋˋ/>�~�Oׯ��}E:u�զ�w����B	�E[3�k�u^��e���IJ��=��A��u����M�AF�x��~�L�l#�K@'��}˟u&o){,��bg. ��1�V����@Ĳ�Gm�a9�[u��ć�K�[*Q��DF���ƶ	}�����U�%@"M�j9��.9;�ռ��||^vV_s�Y4<eeM8�} n���!M[y���e���+܌j(|C�yɼf�.���q6�9C�����沗��c�1F"1U4�wI/끛Tt󴈛V�+����H��B�}s�=$� �/W��`�C=�؅.�b}�Su�$�ŧye�KIƼp,*�C�E�%P]���jeۢu������E`-s$��� d5�=����UUރ�b���)��=ɐ�5��Hf��B�����K��6���W�hKy������d��)`Y�LIMKB�e�I[��G����+����M�����ٶ9�p�F��j��}֪�����u�d��e�{��������7�.���?�����[�V��P�GP��r��6A������Oj�.Ou`ce�do.J�D˝��i8��V��s���.@W�,^I���{�9;Y���N-eɵ}|AMy?	S�Y�$B�Qz�^�%��G|q>H^��Ll@��R`��O!T�����>��W�;HS�W?�.s*����K��Z���r�3��t�j�7�$ǯmEo_�?��@��uğ��ih��C�W���S�e�A�b6��l�UG�G�N��؊��<9���@�ņ'�w�|,Y���W�+Ȼ����
�^\^~�%���>.B��-}���w~�����˻�-7�ύ��g�Z�{�i�7�^Y��~���폗�>��ܽ{�I���#]��_x� ����k/9�N0�9�ur�����/������^>���rG�X|��Um����dk����N]VFsS]42�xJ��7��G��?�+b�q��������מ_^}��兗�W����_\>�����x���/?��O���ˇ��������_t@�A�3��)�'���w?Y~���/o����?^>���r�.O�dkZ�'!���1���a�S]R�
���SSR6KH�?�Q��H��v�4�P�{P�=�5��F�A�,M�պ���y��9Y�'[��kP).a_`1�/�1�P�<��Ӟ����p���9cf�����a�:Yֺ��>I��}��Ha/������tػ}�O�JI@�N��>��=j�'�+��AU�s�xŦ�	p��'�/\��#ڤ0���ܹ3�{(;uQ�3��у�Q�R��G��~�Y~jc#�}�d��o_��"}$ޅ�/�z$k�R��d��{���:h;�S>�!@�&���O��r��J��Ba�E�]����r�Z��}�Ν�K2�sG�����cY؞i>S�M.�&�����K��M��1��%�B֪����_;�N�8ťN��&Tv�i8V���� $�
�R��{�3I��(���z_�y8�	��&�����t�N%h�]uГ*�j�O��bo�ڀm�����d3}�S[짬�d:A/��e�L��R��Z�����!5��[��C�_�!�p;����K��_�'�r|%��l+���4����J�7��l�����b�b��-��5�3&�}�~�,��e?�M^~��y	c�|���o���_�+���nՅ����XD�A��J`rq��C�E8~6� \\��>�&��Zڐ�OP��AP�(�6˲.>� �ԟY�o~�P��=E/�������d� ��=���8T鏯��6���Q�xZ���?�F78�3�����j ^u����	�Q�6-I5�U;��հ�}���7�Jw�)��jw�w-�E��`�?J�r�����]�3ז�_~~��__���ח�}���o�����s�V�S�S7�h*rQ�����.��={syE|_�_xuyE���kח��*Ƚ�ܾ���[R{�Ol�~���ګ/,_�ڛ�W���K_zuy�//�H�
�	��\�,��� �ϴyi>07�X��82�+��Ԩ�
���s�����/Џ���.(�~j��,_����}M�|���_xE��������J<��i؝ۺ	P r���E�}Y������!?����`���]�{�)�p�-��G����[h=da�e�0�<�H=>=�5fd��BG�k0� >p�����ņK�tQp%�A'��|����'8�y?˾���9ĶV��Ϋr�Sn�kos}�e���*c��Ocٻz������*�]����7�}��@�&��G�s�%��S�ӧ5�E��C�1�JW�mn����i\��j.�&�_���k��/����ҋ��=�<���7����r���yh�k=Ï5���M���+�_\^��z^�����p��[�Ƽ���rt�u%�'=���n?P+���L���t�U�k�x-G����%�*A��s�~��Ov%ϯ0�����E�k�Wv�u �T�Yu��iTn�/�W�Db_�e]�E	p�`�b���,����.R�Ctv�2����K��O�G��IP�綺��B>��od���`��]*0<�Y3�R9�����d
�k�s����W� \FV���Na3)YN���8GUy��{A^��Rd���4�*� �:����T!y�Yk��Es�s˛�A,y�@��ȵVRm�!BV�s.�)���>�W2U����Z�7�./��_��ߺ�?��%��C8�QH?��1~��%� wA&�R&Y��2�
pPO˂98*�m�#�͑�j�	-'����6P<y}I	����0"�|��eLQ�}�	�t殊MQ�MohC�}]y��
U�ʿm/-��H?��=���P�>�|m��c���:��=��U㠴Ѱ���]�iGw����ч�:���G2F�g�v&�FR�w9{p���/��|��_R����/>����.��]>e�q�.V�KA1��u1~SA�7����+_zC��K�U]T?������.?�����py晫
�_Z��/-����\���/)0|^��3�����,/��.�7<yϕ�����<��p�簃��+*:�:���r'��@�Ib����;���7_]��K_V`� ��/)Hj�y�6���S
8�R�)	��a=|p��}���˛o���2|
n�PP���O���r��%�ܸvm�zUw�
pϴ�����{r{��Gx  U�EV�(s�q�vn��1��~m�����<���$����-���������Ndx��&"7=�lg�U�;`,�c]���o����?%���OAL�MG�P�y*�X)IQ��� 9<1$ e�6l@g�*�������N���,]?Y��'P�,��.d|^~��_�x}�V_MdU8���n�.>���U��,o~��,����������7tc��_�a��~��[h�ּ~�<��u��W5����/}U/k�5��罎.�x����3>i�MVuI�N�V��'e���yH�`T���y�R�O>(���<���u��np_�^@`��s��5��W��|��u��'���M��~Iu�?������Һ��@��7f<{��_�����o>uSxCA�5��旛,�������1����]_u>Y���!x!F��o��@=k�	�l�X�g�~O��}���w�\�5�����uZ����C6a�|L�����B�_���峮Ax��U�c�v�g����1Mu�<m����I���xΧ�A��-�C�d�m�Qu�4�W�T�/)��$�1��-�'oߊ��^e����8�e�	,����~���L˦_�1�<k����M*��Kp����������B�X8Q1�B���xp�DM2UXV��7���1�cܖa��T��$,T���zZ;R���/z��[�G9#OmM(��#��Z]����6�\��T��Z���Uj��9�Z����F���^��N�M�ct����Q=�y��s�3_��i�}���7�UǓ��C�+���Ǚ�Ǐ9�����r��^��SWؾ�|�<�|}����-�)�v�'$���\�z��1�����{=��B�ګ/)�{C���˳���������w�}oy�?Yn���O�x:��_���Z]���
_�v�@�L]�J0yC�٭ Vr��UP� �O�4���'�'x��M�＆�k.�=�\Pۃ���3A���\_�� �K_�	����?���.�ǟ|���r	s��T��ٽ;
�/,/�B��^v`��.�ׯI��۟��}��rI:/��{��5���r��O�,�||g�w�w�3o���/�)�?5�LJ1�&y�BWD��F���!���i�qˋU��NB�8��w��W�3p���)���y��9N������Ԓ4�}��F61�_��*r�o��`��;�4�m�/��>Y?_�C<�jg\�ov��G��u�O(�&��#�B�P�+�Ø�>��-�CW7�LO�D�u���3�,^^^y�OK�j���S��_QP���g�g��|���<�<����E7�O�S�_��ٛ˗�ȧ���6�L§<ݖq��|��L���������ut���{�l���m~����nyO�D�o�j�_y�E��//�&���<���:_U �}o�����k/+����+���~U����}����}V7�������n�q]�����{s��oq�mg�3��zʍ�5�{X P�>�T�T�1��&cR� �>����qG�EX5G��i���i�}]g_�;��,�|�Ķ���n��Ÿ�k�f.$>	�}�wX|:Y�*�(��%tk} }�kL�k���qƜu^}G�`��\�)?�K�? ���f
lg��N����%F���Q9�X�j�aG_��������9
&E�+�i�+���N˅o�ſ������Q��2B�a�lZR�'l��,(���/$�U9|B���!������JN�شwXC�GήI���	;x�b��w���v�IR���>�J��<�E���b�Ƈ
�%�@��lh�p���b�ye�DU�}@�R��D2�?�R{�K2�������Q�a_n��M;Rr|~(�	Ƽ�[�+��.��穀wO�H}��_\����u�|ay���\�=Z>���r��`d�b�����y����/����Rp~�����{.o�����~�{����o8�����U�_��ڋK�'��ݒ���<�)�7����ɭ;
��-w��_�+�up����"��ugy�$���i\���Ǻp���m�@6+@���կ��
(����3��ѣs�;�~�|���|�{?^���'˝[\��R�	�����������ڋ�o}����[o-����,?S="���`^A�l��;�G��I���:^ޱXs�<m(�z��*1xc�̈/�d������'��u�~�YAm_�<��{ؤ+��E�2�o���m|����%>�	������d�fϾ%�<�'X�SZ�hs���h�3�H����yǔ'�޿D��aEʡG=>O{/������'p���'����q{p�v�腍�)�.$J��.� ;My^9�z��T>�=܌qc�L�?~�������o|I��ۗ��}j�~㊂p��]��<��%��?��������A�_���i��_���eݘ������K�r'k�����<�Ⱦ�@���ۺ�R�k��Yk3�)�\��Щ|����?sy㋯�F�k~j���~Q���o����������<���K�[�|(M���g�7�������7uc��s������v��;��5�tzS����������_�n��4~r۟���E�~pʘ���`$�q��L���t04yO�k��f�d��#��^+MoT��uY�ڨyK9��&���0�(��F�u�5՟iM��� {t��	t{ˍ�G�LO�p��LWk�%�D�����Kh�@�w>��T��Ū���G򴶉�{��:�e�Q%s����u�l�~�A��A�l�&��F�*�On������_����;�H� �e�7
0rA`��'��������V<q�������1!	n�d̤��������l7�
P��x��()+�	q^H���oL�}������[(`<$]���*J iЛ)H�EDN��?磴Bц�x:�Í:uʙ�S�*���� q�a�"��@Rhl"s
t����p��| ���C��aq�?}x��]�,W��[^~�嗾���+_~uy��E�p����[��{�,?�����~���@�害�����m�	�x���민��u��-���Y�z���G?yk��?��r����W�S@���k��~�����'���������/�]Յ�_�#M�ջ�}�|��-�\�y�T_J�u'92j>y<�L���	b���E�G��_\^x�Y��.��,/���l>�|��������w~����}��?�����ꯂ�۟���	/�����}ṛ�����WP���'?��/�W._�G�|��4x�緗���d���}��>��/���N�9�E�?��e�M}���A�_�5 ]6��F��&��D��+ʐ��ru��k���V~�[����b�8��B�;����z�d��l�΁H�c�ai{���_{+b�	��Q�@�f�����%�?�����,�`�\���|�͒bKA<��*�>���~���YS��_d�}���"]��^<�����k/,���_]��u��^Tpz�7b�uC��Ƿ����O��k7�sc��o������/oj-=��Q^C�wW7��|��������%ٺ�Sr�f?��c�?�&h^����o�q���oA��c�~�Om_{����_yÁ-��Z<e��B�>+�y]��:K��޹�ϯ���򕯼���7�*� k1/~���Zs-�|������W�����Ez�$��M)�E�ix���nc��,)�W�3�y֌e����x>G�ʮ*��v��=�fz&�*�=�u���w��(ٶV�I�J�:_4NYG���[p�Q�[啯�A�V�S�i��ӆ��4p���*�|�-������f������C�ʠ��.��W) �{�j\��#K.��භ ;ۙ��Hj@���R�VR2-k ��%B@���έ�k~-����[wt��O���)�Sj l �"��"K��2
k2�ʲ�$L@04а�c}���
D�S"���\:+�Ğ��VU�� �o'�	Oe�0���f�51���Ke�:�K������
��j\q��J��6NiSj���,�R^�E�/��?��z�l���.��rR1�`lZ�#(t#���VI�����@���kE -:'s�~���9�2
�W�N��h����|B��B�nˇ|���?���/ey㍗t��������/g���������?]��-o������+�}���=]X�=���D|�Y��@񱂼����Ͼ�#��ݽ��/��|��T��e�;��{/���]�����o���.?�����7�zn�y㦟@�S���[�K������m���o��x�'����7=��t���A��fu�}�g�/}�5	�i��'�?��O�?��?Y~����{����|�|�ޭ�#��+0�⋊�_zyy��gu��ԙ��~�|��'Z�벝'lO=sC�^䷏�( ~O4��3~�D�(�:�h�6P�ެ\v߄��ā����./c.�1׃��fQ����؂9���p>����9�M ���i�2�ϛ������9������).(y��6/�T"S���a5�����B[�',��٫�����������r��-�m�w46�����j��^O����N��{G<w5��6�_��u]�?R��sO�l.��0e����_��������~]�+^w�u���T7�?�ty�]��xI��r�S�}��S˫���y��o�߽�O~���h�Hk�#]خ�v~��׈;�����皯w�ܓt������,�@�[��ǌ*Ƒ'����Ӛ��/�~��o�U
~-��@���ua=�h�-W��W�Ȗ��	�(�د|�'�/j-��Z��~������������G�ȶE����__�ܯ~c���^�M����?/�+>o����ɫ	�o�_���	9͗Tsȇl��)ig��)�eH���OH=�d�n=�����+�7�����Z�QZ�f�e�,e���sP�XF��D@2���R�D,м�qR�����������U*1��2&�1R�H��C�~'m}e#<��Nyw�\tJ���)=�ϼO2�<�E���_o��v���.tDU���A�����)��Eg1��-(=�'J�e��ȧC�)��|u�J�
= R��ɀ�R�"��!��۰=���&�F�<�=9��2�v\���h�7����v��M
2��.b�)�C��Y�ŲA*�PF�SՓvP�����y���0ߜU_Dm�8�	l���,�^�5�6C�����npZ�b��&��h��8}�a?B'�1���`Ca�����u������m���3�o�;���֭������G�g˷�X��,d����_���-?�1?	�����VPJЖi�5t����@:&.]��\���G�t���O�[��O�Lz��|�;?\~��w��`A.׀�;�,Ћcc�_�A�I)�^��5?�,h�11��@x�R����P��~��P������'������?����'˟|��ˏ~��_�8��t��\�~����ʫ
�_Y�}橅o��~'������|Ҷj��h�1b>�`L�=T�YxƔ=���Q"S�D��u׆�����A�fC������_�+:�a;�|�~|>&�Sr�W�	hA���N�!#�ӗ�o ��_F���2�:���^5�
h��Ś�}��������9{tG��+Y��(P�x��͇[�r_rry��+3����w��c~"랴�4�/A)(V_���"��s�ϼQ�'�<�}����O]_.i�X�'?~{�c͵���?Z~�w�H�x~_ﻚ��P^�rU<O��Eًo}|�s�goi]���/��W��ƴ�6_��Y��~fM�|QE����aT�}�������5����U�|���M�O���?���wtC����
p�ǧ�Q ������k
��u�g����_T?..7�]��"�@��ӗ��Ћ/<����S��ϪϢ����'Rܨj �(^���T�0:8��:A�Mϫ-X4��c�������r��1bc�z��3y�"�(�jα��"�Aץ-���=����@֗Sڴ.�:�ǩ=����h�|ׯm+�uȩ|�j������H�C��9n���^�6�B������8��2��t{�S�ed]4@���0����=>�3'=^u��nkt~�\��Xδ藬��A�?XДZ��)�иB���_a'b��i;:_�h�=&�3
){q�m�/��^LԞ���!UZ�m��	v؇�b̷�٤`��� ��`��.����I���v�1ע�O���?ۇ����9 [�v#�R�`@���dr�y�o4W늾0�P�~��?�	���?O�����߃]t���~�@ݣ�
R�����������~��?��o;�㟼������B�0��_�c$�`?���x�1���.]��tq�r��.���-�^s��WXS��UY���S��n�7	)�,��|� ��-9�J��@��-��.+�"�9�����
������}o��[o-|��r���r���e]���K_[~�/����+���/ű�����=��s��0�ѝb�����62�!�vҀ�Ɠ�-����P�"�lI *Wh̰��;�<�|���<�$��+��'�'h�=n���o��� �c�|�I��N���w�_��u#C��Lo��BT.s�UL8�/}d�k�'����
���`���t��r��'"?�nl�=T����]��LRtӦ`��j�oi���u���W��W F*��?2�7��7e�|���7����ؿ��a~*+{O�����~�;�[����d������_�����_�?������`����ǲ�CIy`;4u��n0���Z��߻wG�~<�oX�s]��<nP�:�o"Doo�?���2{\֔�׉�s����ʵ��=�����������׿������.���������) _A�]�O�B���.X�\���Z���1�C"�_ 5�Ga7X������W��9����������Eh�e�'AGɤ����oz���_/F?9ʾ�.`���:�\�����A�8u��1�7v��.K/s�X4+���k8�g��$�<w���=�3e���B��f�mp��4Ӹ�*L )��[R9�:R7�I'���lѢ���Y��ka��*�~M�a� 勎�>?��'�p¾�� �vGG'N�$J]��Y���HY��rw�uVX�v;G�j��1W��L46M��	�Q��#�oW(��S�LH[�w��cbMX7sT�h����8��XS�]a-t/���; ���K'&;f*]��y��a�3�3z��olo�mK�����&A����?z^�������IO��I�[�>Y������o����ӷ�裏�e�|���z�c 3@̿�����Ȅ��r��R�9_�z��Fδ �7fӍƴď�Z��Q��IY���J��?�U?I$��	.���7�yO񲢔�W���痳�g����n}�|�ɇ�'w>^n߿�����חg�{nyᥗ�_~iy����(��`��v�7��s���.Pޝ�Ƨ;[=>D`��@]�z6��+�Ws�~.��i��!��G
��=�w�>�O���w.0�!n`��O� �A��Z�<T`l�,�M�"Am�L����e�_�@��#�P^���3�<�UpwN���2%?�o��K�]篿�|]�/��˯��?渢��Xs��r���go����8��xs��o|q�������_��k~��Ko����î]���:fW�n����=Dv�g��qcx���ˇ|�|��0���������?�S�L~�����G?�ܺuK�W'�/.�'A~U��W_���M�`��2�3��������|N���o7:�b�+��f�)䎄���Bp��{-��?���,��;� �O����?[��G?\��ݷ����go��|�����$���lZ�0z��߰7�њ�u�#�4���O���g��b��fL;����]q���5;�NE�o�'��~�f
nh�1��[s}��_�F��g�ޣ�b�:9�}eR�ۈ�M>��h��t���]|��H�v�~����糯��������Zm��i�C�4ѫE�
lh}s�ɀ�>ZL��ԑ�έ�k�(�DqW;��3)~F�(�s}c��[�ȧ�-=@M[�>��gˌ��8�WTezv�v�O�)��|�H"9�H���Ȩ���yOX�*~�'e�0T���0�T]h=�U?��M�������`ߙz�@X���>�,�b��,8�7wO�`�]^��3f�qG�g����3��^|l_����ɧc��&��D���+�GǏ�X�'���d��=>��'��mj~W��V|���嫺�^���4���P�_F��<wA_��^5��4&_�:�ϸ�-N�S3�P�8e��3A5���GҺ�D	y"�?�觉��E��h	�6q������n,Ͻ����+�,Ͼ��r��x]�/ɶ�����������= u[om�D!�.��`{��{��~����2t\ ��Y���[QZu��g��)�p9�S��4Vh�>����ܽ':�F�HPk�_2�6���r:�x��[B��tKװ;�WPv��Cd�It���/����k��
�;����E딧��dk�$;�!���+�k���|�W����������m���������󷗿�w�����;}��_���������^S�����7���u��//�o�����o.���W���7����������7���W~c��_���K_|ÿp৔��c/hL@�R��E\�uA��n�?�]�����֎��n|���ˏ~����?�����x��[o畠�n˧�����+�7�k�_�������ʯ���G~:|��k!{C|-sC�1Ә:��g�!sFk�!�XHХK�����c�G
`��-���������o}{����-����^~����_���/�����D2� �+A��ﾳ����������(���:� 9�����o���2��En���*��d\?J[��m�σ�ܭ����sr�Q�,�%v�G���C��u`��yr�k��6]���f*m�\���Q/��Ͼh;r���%3:c����d���JW�3u�P���7�[����
?�Nv0g�_����_ʘ�k��-l�+�>�I3�e�e���[�!M�`�1��I�#k`��.���F:)�S� �m�M�ts����cțe��;��+i�d�8 L5��]���A��L�Oi_�6Ȇt,/������(?-fA�b���cbr��b���S�t�%��Y'1��R2�$�m��Ǻ�݋�4V�I����?�4I�4]L#��ΓD����}n_\� p�s�����+��� �� ˙���=���3#��s�Y��������ʪ����j�DTDTTUTMM-��d�W	�&�u'K�e�����g��#�k�"A���w�{dy	�}�c���޸y����\V�X�<�(�u�� �O��B9�k��R��Ӝq��W��j�"f�0뻠��ƀ�d~��u�,�[1��(yxp���*��-�O��ə�6wm����n����ۃ�[�n*��b<�z����旖��gOۓg����Z��aO'����Y��;� *]1 0B��W�}�1ߋ�.C^�9�W�d���6T�e�v��}�ԥ�v��T�)����������ߕW�S��:{i*���c�H�y�/C�5���y����[���������+2�d��b���1\��_�{��@΢-�}�J%�����킌7���2~�^���۟�������~��/��������g�?�����|�Gvݺq���ه��i���>w>���4�g?�L�i��s^μ#�xN�-m@td��@k}���;\��@�2�ݩ"���Z���(}���S�Od����{�U/�����܅���~�ɐ�r��,IK:"1�ʠ�1�6�S�����%C{cm���m�Օ��0�ܞ?�o�|�}��o_���<Q8��&Na�Fi�^7OԮ�7���B[^Y�����) �)�m��[џC�����r؝�ǝf'���f����"O��/�Y��ኖ��A�t�m��@Ÿ���H`?�f���kC���2,����?�}
��
q�a,��{C��}��7zʔ�[fLt;�U;(����F��d�m �Y�tŕ��/GT^v���q��࿜y�n�PaC��y�>mE|��Đ(\Yf���{�sZ(6=��
��{A�9�w)+�|9Q��U�PY�]�d���]>�����n(1��4�p��0f�Q�D8k��'M��־:�2��Mk�V�x��3s�V�<�0z�'f�qm�xA4(!���[@�j,�F�Z�5�9�n�'7�HW,�Qo�&�Y≮Rz��ċ=�#�9��xU:�&ifU=���=א���+2>8����	�(p��e6wڗ?�����?m?��ڇ��K-�oo_�//�`4��zԄ�U�Z�
bqH;FU=��15/�p4W`pJ�d MKPɳ]dl]�q�S��z�0�B��Eyk{�(_���������_��g�g��Y��G_��׮^�n#b��|����w�i���u����ߴ���k�(��t,�������7��B&�@����y	uo���Jw|�0�9�LFb���Hٳ��Qn��&m���ˏ�/�e����e�o�����������w��ߵ���_�O?{��O�P5�� ���x�!�<��,�bu�ڴ?�ˈ��Oۯ���^Y|��ߞǸ�]���^R�~Y�"�̝�ړu�{�����#�
}|z���3�~�+W/�@��Oڏ���}�����7���e�ޝk��\jx���/?����O�s�f�~M�:�7�n����c>��{w}�'ޮ�@��& 2�9k�M�r��K1n��e<>�g�R7Y��Q7<a�6md�Ҵ_����p���������ۿ��j��~�~��G��G��W����/��[����Z���	"*/�᝾$t}��.Aϕ�1�.���Kp�O�9!�D*���2�8<o�?n/�>m+�����=��́�k�M����Ͷ����V�ۦzNR�Xܦ�?�i�"eH(<+�ڏK��0�q��/0�����_N��<\���]ׁ�u���cI��j#�a˘���"t�A �t=��*r��3I�L�t=8�6H '���h�����=Ы��}��>���v+P�� X�@O搝a06���[���4�uZé��ʋ�(���6=D�5���/�K��e��o�
����Gc���.���-��"��N�x���6���P���ua�#�<a��x�D�$��*��١*pwe�#HyQ����犂&UZ5N^��#��z`g���eh��=v�v���a�����Ip��- 82m���4��q, ?_�S�B���3�-y���F8#�Q�U����_��#��3�!����������x�?�4N$W����K�t��;F�B.���S�v�`��^[����!�&��k�&��q`�����g⾯��֝�^��`|u������*��G��T&m��>qx��s�����2������޽n�jl"�Y^dceH�hp�:�$����H��=U��5�I��ș��Z�&6�|�"��x��'��/���?�P�П5}�ч�Ν�mf���	�a�� y#<\�
�S1rL"X��N {hHن��q�+C�q�ت`�4}�U�Z����
J G)��;��o|4ܭ�׼�������|�~
����������ԏ��ҍ[w���K��G�+�JpQ�._���	чܓ!����g��_�����ˠ�^�7tvv�+��ׯs6���ܠ4. �OY�o�q�G��~JA�k�8��ԫ�'m�n�@}���ޗz��6��<98nj''mL�u�꜌���h:�D�8�c���������fwp���o��̔�˞��3Ӓ�d-�Ne��/�V�y쉑�
�P�gr�1��Xe~��n���[�A�-�z�	�d�+:V�7ۋW��_?n���5��c{��ElY@�R�0椇�ŋ��t*}|�pA�/=}�1��=(� �RdO�S�hKx�63,=B��������|D����Xn�{�NK���+�zc���e���qw��s�=i&�\�mh
(Z�"���6��ke�l"M7&$З�Q;n�Y��wc����d�,R�a��^�k���[i
G:����QO�� �Y��C�GL�9��r���xF����2�ϧ=C\���q>�����ׅӗ��@#<@���N�t��t	x��p���gL$�QƾA_�"�4��:�#M�'��˂qD@.p�u�su'ފ��=3��9��*$���#���r#��o����'a��LM ?_'1n4�Q�Z��Rp���cq�`pAY�	%6>�dC�C~U��Q4f��m�}���u3���cOMt<�/f/�T�őFC!��W2�N�̆ľ0dݟ��~V�H.I
�4꠬�4F�vb��e�	�H;�a����� �&8\�9�W��Z��ٿd�� ���~:�"�(�0�E^�LCz��}��A���wפ��y�hhsϵW�|��Pu(�����5�+�D��U: ��#�AA�	�W�qN�`�MML���vM����ۇ�m�����v��6���@ǉ�����ݻ)_�����F�:l++����́�e?�����/M�J�����I^�?�+D��fmm�=z��^ͯ����9
�ŀ�Kx5�8¸�81+�0��e8���i�Q�2}��1Bf�E�D�zm�ݻW��/?�w�o����R�T'�;�Q`x��8'��&~޻_���/*a،ɰ��=�[mqa�-/mh!�1H��>`�>V���P��Zq��]+�Ų�F�VE�b��5l���G%���:��C+���/R}��n����U��t�QLssS��	�l�븡��ӎ������!CoW������|�����>k_�H���{���o�[�$�i�ۇmsc�/��N
������ ^��s���s�Q|�]��~yM���s��O?�߻w�]V�c��/�'_�l�/��޶��c�gTF�Q[X��Dxi�@�����S4����%��yʫ�*Lrx��7����N{��D��S���k���IM��J_� �x����Kd[;[����kx�P�~��cM H׮��	w����Z��|pp؞>ޞ<{���=)�y��銍�ã�mm��--lIW��恪[�:�`A�O�6teԎ]��m�-[�'�?Q�ЎTO�ի���A^`��Y_�h_˸�S��F;�ruF��+��;�㼵�.[��T�o��P�|���^I����^�?��[���]���wo�{�I�K�jCK�k�����4qe�[��YC'�]@hM�� �tW�y�b��x���0GR]���;�W���L���(��1B.�:�!�A�ˤU^�m	�פ!��p��߈"!̧�:� 9N�K����L/~�Ώ8R;e�6�eT��ŧO8|�8];{���ZE�\�NNۯ��!�����J����5�_"Ʉ���V�n���t#��属 �剕d��{�Q}�}2F�ł[ȯl�2�ꕟ󉦑q��ob��p�N��.���ch�|2{By/kl�ʭ��"�F�.�R q&0[�
��D$d���*3=���{]����.q�D��]�q�NX1��q=L�*���\���O���T� �N��B!#.J֏��Gz+k���y�Y���O��8Cd#���	@'���b��m1)	%��Ǆ��9_P浮*,}@�|�D��t]��V5
��^`����Y���-](�W�>�侌��~���viv��e�wbr\����	��cWÝ����|��^����WH���ZG1�c�b4���_�/��D�=�2M��{mqy��m����tТ?�RZ(f5��,�����f�����Ã㶱���q�mnq�7ni���C�����{L9O��x�g�g��+������Y�ex|�>�q{��u�aB��ͮ_���`^��ژ�]�1��+���4:�¨��t�u�a����G�Kq�?)!Y�V?�Ѝ�+��Jی�W����nεK3Mժ$��*xrT���_�D��)�/[I�^�@�Տ?~��>�c���J.g���r�?��TzP/�&�*w�øjk����/�1�3|$�Jbn[�5+�2�/_�iW�fڬ�����i/�-����W����o��w�k���G�?�j�6dxɨ=�q��c�~��?���i���ߵ��~"�w�m��{�5LGod���#�؞�^QV3Ec��c-/����'����%����q�܏�E���$����t��O����nJG�j2u��M]ߒ�|�]�u��ʐ��e�ƞ��R�1�2��vOe�z�qO���Z�kC��^�g���4����G����͓.O����ҟ���n���~��'�O5Qz�Y���7�צ��I�E�̗	'�t�S�O����$X�Ȱ���	���џ����������V�c���4��oO��$�[];��b��1��+�e���0� ƍ;��$��*u�Ee$P<1�#�7�Y������W�o�,�����m��tf����g#r�U!�
� ��I�FK2��ք�_��y2��_%t��_�/�1ɸ,��r�[��!���
�<_�}(y�s�;ߘ�̎_P�T�+G���3����2���˷A��7�������蠰m*��`�����Z�H�����U[�����EOlQ +�(�����*#+"�����Wg��C�H��'��0Vn��/ �q��|�(L�y�L�5\��7�=6�����g�����.��L%�r��BTfB�;���V��.�p����ϵG�!�����_�"��ex������v���W��L~�0v0T��2S�]�3���IKD[:��"�W��� Ʃi�A:55�AcZF���h�������nm}�-̯��/d��I�I�&��pnnֆﱌ���2L���ʚ�CO쳝V�~�ʣ\V�yو��!~r2"��=~�*�R�c����SRQ�B��F��h��I�/:5�Ι�n�����)]Ʊ_�4Ƕ�q����1��+ߡ�������h���������acgdl\�)�'x�m�DDnn*�F{�x�=}��VeLo���uO$�s]X
�`��G�W����VE�ڵ��@il��,eᕂ��-��S|v�+�_|�q{(C���e􍌢ݶ�����zۑ�4:[M$2?2�XKKK�2'^�i��_�G��O4!��U_������۫���ٳE�"��Z'��bGG'�LL��O��;��'�0���"���xi�Ht�7�����۝�W�ud�5;����o�n������^p���鬮m��ն���O,/q�"��$�ޔN_�$�v�}�V��6'Z��FivT���q�-.,���}���q�a��w鲌Q�!����x��4�n�H|���m�>�X���	�&e�>�6��ם{�4!�"�ۇ?n�|����y\ڙ�Ot���x[Zo{{�CO$�	^x�ie�)�}���(�	R�g������׽���y�¸���z��'~�˟hr󉷀��k>*A{�%C����s��W�io{{Gmiy�mn�����D�P��o{���/�GlǸu�O�^� ���4�M룺$�9>��
�_�V�!_m�#�]A޻��];"�y�x'd+oP�p��4&w~���ۑ����8���t��d���W:&��x�jK�6b���3�>9D�9<r��C��t����r�;=�u))��(#&�nO�������GF�Ѡ�1/��«�ЗH�~�*����&����=���Y���j�����a� s�^ʞ��geG2)v(�^�a�i��xI�v{Qm�'�|e�g���N��q���=g�a2V�@ �L#� ��<d���!$�[H��	���G$	Wr��_ބ_�:cT i).�4*��@�7n�Ÿ
!�-|1���p��ׁ�\&�a�I\�g��CavA�]E�:o�:�
q� q9w���9(ʫ g��:���O�	�_������]���������"���S�o°t&�ǿ�g��IS!�x�)r4&^���&VDx�>��}�O���U�1'�+�ϟ/0L�����I�-��A��@���Q[�Q�'vWV�e�h�:�2 �tM�:NK�0>��wҖW���}����W�k2�vE��M�0~�`$3�Yi+H.|�LY�{b��c8��1�^;:~m�B�+�KK�2�7��_���z�$#u�o���0��Cʷ�w(�氭o���-Ѿ*Ö�i�۪�]�s*C�@��4X��-�$��ʠ ��\�~�7:�p(��mG��ի���&[d�chٸ�{�}���^e����P��W��=}՞|�\FҪW�ų�������bM�=�Ӈ��Kx�wnߐ~�~_Fժ��G_?o��T/���J�*��B'8#��N��`)y�������K��;�<���}����7��۽�7ۭ��3����[n��~�~�/��;�|�dO<nnm���-�ߖ�����^�=�kC�Ա�)�Ω�~�=}��s__���t3:B��3�^u	]���{ly�R�=�&_�kW�]���65R�H=��&��;�AF�&!��;w��
l��a�8�d�T:�1]�'�!'�E�#�#�
�@v+��;�2n/�btO��A_M�U�ɑ��l+�,&��0����ܼ���dp� ����z�@u����;|i����hׄv]���۩�	��������?hW����iDm��hG��p��z]�o]@GRw�S 
�y��&�ſ�k֭u|�wO.��3�����W�ꋥ6�z��i�䓇��F�h�6Lu��n#V}�[�	�o����q���d܋.������}�=q�N�U�Ëv_��e�جB����1r����?�3�y��4�Qg1	��p�qk?q{�D�x'�a�urN�vu�q�"��3/8�G8Ҏ�^���&.�����F۳>*��m�c$�qw�q������4n�3���ƒ(S��!VNF�r�ag,�r��)�q�V���I��_7v���[�$u�e�)����T5���S�v�)|(�+/�^�H�u \�.H)��'̑�$_���ׅ����g/�p����"H�$��G/�]y�Og�%�>Ic�U�`KNg9$���o9*.�v%��|��𜔔��W��$"��s'\��"�\�@e�8�E�1U�9��W���<��{�؎y���Z��kk2T5�,.2l���E{�t^���V����h�}-�tg�Di�N �a�6��������}����n�x�#�x��B��}��m����l�<^���}#�����U
ZQ�N!g襮J���+����Q%FK�SG���6	�d����t;�iK��f{!����+2d��`eyӫK�T�og_��*�v[Z�v�gʋq�L����m�-��A!rcEF�d}Z� �_���tyA�!ׅ�BP�+�p##]Y{i[2�xL��������n�S�2F���>��nޜS�~���>j���߷��ߩ�����+6L1��={.2rXa���~,�cY���j]��Ǐ_�������?�S����?����k�Ϟ��0��� ����p�փ3�=��/�O� F+�$ɕ/�Ez�g�Y����lwD׍ks�%��IG0p?��-:�h��M����	ܞ�t_�wd���������?o?����'����ݜߦ��V��^���_P�� ���o{��ˊ[�(
m�z(����I@�P6���b�z�#��������6r��΋a��Wڔ�\>J19l��4�ۓ..:߳'/��
m�}��'��'ԍ{|��cɐ3�����ls��)�W�/_��f$��2�gfgDǘ���sҟ�ޮ��l�X��`K2BO�'Wۭ���]�8]�B����I[�`b�+W4��k��4Q��G�iBr�ŧ�����mlj�w�I�d)b�� q@����.n�ѴA�ȧM�=\[�p$�Ԋ|�a9�x+�-\�Y�b�'��t�)�������~͓t������2b����X�(��r�½�T�p��jPF����L����9O/��ua�$��_ ��Kڜ���WG;?�6����m0/��k�q7�)b�O�{Y7$�a[(@>�'�PWG�􁇔,|���= �mK��vĻ����mD���0nm��7�4�
@ق@�pA�� rA2ƈ�N��}��HlK@�J�@W��1\���C��z��H��|��!�>u.&�IP��G�SE:�#C@��J��a:q�
ŏ�����v���<�'�xE!�tN�C�8�ɝF�e)��G��A���9���r�3�����rʸɘ�Oa�θ�0��]�&��81u����"��sn�ʇǛ�2�v�5جﵕnK�maaͫ���1�no�9V��Y�2���V�do�y�+����@�'hc �����ȋE���/���/�5�˸\nK�mS�cآz���v�AGo�,��ڠ�	�r��"-�^l%�~��˺hX��r_�(}�L��+��}U<q�'�C�'Lj�1��2�(~_�Zm/�-�y�_Y�i�k�m{s�m�ߖ��1}�y��.۱L�q�-'>�:+�pIn6�D��A/dp��Ő��۷���?�߮�`Ae8���Ծ�Q���3��[�mkS��\]]����؈����ۧ�~lcdf����J��j�X��Q,kS80�'S��s^��u[t}��+�Af�Ī-za�6�*�r�d�6MeԎO��K����>����K�/W��/_,���>�R�����&<u@vl`�'�~�~��/g���֑&Iϟ�R�|����s�<�wt�=���Ɗ4OK|���?�Zz(;����<�@ƞ4i���劌Z>g�BmcA:����<�4ϜF���$�0[^<_�a��YȞ��1��:,�l��0ne��C'�3���QN=���t`x�V�1�}��:����R�9��-Z�Ԟ4	�Ig����j2p�[��������@�h������U�wn�{��*ό��;�~�W���]b�3p�����'���~�C�G9}�G˂+�@�j �y��wFV��х����~G�#�`��Fхs-�G��}z\�-�����̔�w^�k�u�]�A[&�.�����Ti@lǵ�3?;�;cFAj����U �(l⨼�8�_o�V�#'C�!d��` /i?	�8�b��޹r�$�I�!��������&�Iu�|��!�p���$�:rƸ��_и�dAU^�)
싘�!		|���<�� ��F�q���b8Vn1n�.��&7(oK �3�Y��������V��O�#K_In_af=i"���}�wT���^����K?��L�&�?��t���BII��D9�{<��뷜�	pp��o�t��#�4]�G:w[ _�����t����XyWt,*(.��x�� }�|tm�mU[�l��X���{�}.��3 s���چ�Uf�2TW����c<�gP�)RKT�Xo=��va�G���rѫ�*k�G�;*�D��3�V �e�,$���`W�8F
 ���6���8���7�y̾��'�4�.�������j�-/�)l��A��=�����G"nw���7�v�-��W2<��˚���V���[�w�'�����C��s���N��=�|���O$"\�O_b�!Kw��؋�ُz�����7�����Kt��X�jOdTQ/�2<�v|�){>��6��y|tdC���>����׽��F��au��~y܎Q35}I屷Z�v(![v��b�Bq�p�w��,Ot#�J{'ֺ�+d
�6n2�9����������^�B��?}پ�����-�ek�3��4fC�:`����[�/>�^ҏ?��6��.z�o~�X��퉌�5����C_0jK��:���2{�9�������˗���G/e,���oT��y�zX�1N=����,&f����ٓ��B{���x����m��o�� ��R�}0q�_�=F�#��ā/��n���Yu�%I����'{�/J7ި�8nk��.h��v�g�/�}���~26>%.h�$�vu_���yɍ	��+�33�D�?]��`�бx��	*˚|!3ڨ_"oq|�X���~���᲍	���Hr\�����n�*.⇢T�Xo�n�q[���U`�YG�V=�i���?Q�[��q� ���ːԫ�x�*�쁍$���oi�~�>
�-���H��S6�r�H����Կ�g|��k�o9FoK����g�M#���y3��OZC�u"��	�֎,�[#���zz�a�Vrv�tܻ�t�f�#��F~�w�����Oer�h=<�q*�gd49
����BBH@0�a����m�zF!#�{Eظu# ���J<ര1f �U!�p��6n�t��\���?��ӽ���^�`'��G�NP� ]�s�/*x8>a���Ɵ���e?��|o;�'��qw�xP�z~Gt�S�q/�3<�2T�~y]���X"{��n�4D�������K�hPg�$�H.�"*]C�r�({!Y��E���]��Ǉ���]�4���Q�W�4@o)�
/�H�E��;�c���mmrb�����\�v�7�1X�S'�.1{e�e�����0=������n��?�SzV���/�2[$d$��#�t��?���7��+㋼�?�lO8�ʷo~����8�?ahb ��PK�B���n�D��!�z�����K�(����2�~�֦��ڍ�W���� oc}S��3U��{2�8������''��~�񗟵>|/
���9��b�>;;��iΌ�q�[��޲�ʿ?Ӭ�1[ԛy9�<I��c@>��ҵ���m�q{�]VG��n��e�3i_ZZ3O�>���}�<j�}�WA��nܺn�����Ï���.۰�_�n�ͷ������+�VY��S�=`��~��6����y_�6[dV�5��DkQ��Ͷ�I3m�֫�V|�0�$k}W��v[ZФT������9�0&c�%r,�0�22�61��y2�l���"}~�ʭ�-�3�M�Ԗ�N��ƾ�SѰ�.C{MF�R��3)�d�&��϶���}��<	�~]:Ǆ�z���_p��`x����6�/xc�1gV3�4C8X�2X��e��q�/�V���]w�2�l����ez;}^׋��=ȶ���v�p�XH�"��,�vO��1�s��X���t5y*W��[��
LSR7:��Ɵ�@�x�޾���Q`�1n���?R����c�|��-r��0�#��W|��+C	JF�k���*6�"�#{�y:݇q�����x�` a�(.+.*��tO%� \���NA�����'A4P�� ���(�������u�x��Ap�Q���%/�)8d��0R3��Bǆ�/���" (��+Q�jk����)<��f2�A��/�[�3�0d\Ɖ]�S�m�si���)E�]>H0�~�������{�w���/�k��,��~֑��Y1t�o�G���S8�>�:Z�[4�QGX��i	������\�x��3.�z�� ��tR����ToΣ��	��h�8�t�4�@� ����yr�������x�,nVQ1p��X�+�<~�����IU����Q^H�.#�_���U���)���C}X@hl��_���>��]�9�j"�=VD2*l4����j(������ĄW��'�e����9{ף�� ��8�7�''��O;�
QY��>&�Q�no��hwvuin`�~�}/��/P���|��q���ХQ�餾��S<�b����+���*��GO�Hys��hZV|��4�8c�ڍk��ߓ��Y�'�����uc���@vynʧp��Č�Z���+�词�~W�	%��s+�5�k�h�`ܺs�5O.8C=/��]�i�ߕq{�]�2k^X��������ȧܻ�}��/���HF���s탏�k�~���}��������q���e�>})�(Nݐ�J��t�&�����Bo�;�bЎ�����zh#w�ɖ�^&[� ���~�(2>�~�Q��M�v5�ae��dD��#�a�s�	��\�Z�C���/�\��!����:90j'��&��M챇���˗��]f넷O���b�OC0zنē��}������������z�"]ٕ�⁾�6>����+�vU�����zϷ`eeÆ�����ϴàB�9sz��������#]��p����Z���k�H��� �?�>�~�ڥ��?x1��缅#6
�F�x��e#K�T��F b�`�}�!�:!=�S��Ls*�KW��y\'Q/�� ��y��Mn�w\��@^ll,�+,8D������9���9�-@z�h������qe����F���D�B��E+>H�%=q xE�i�X�'�t�Exh����%V�u_�8�A��.y�<i�cۥ��0n�ԉ��|&�Ȝ?�2T'�F������B[x�#
g<9��q�{:m�y#��;�ș>.�Px��pr�a�b�&QA�խ�"���=Wq���h���/���Xi���&.� \�e�{��p9A�\\�%D��1�v��W�	��__ʝ�w��W���ví�rd)�$Kw&e/�H�4p�T��0�8-�-���?�C"��QxM�.���`JS����HSC�c�����ݠ=
�����#&�y�W�D��MMP��n��3��ȗ�4x�N�}��%�J�ق�?�����I�iȸ���r`�J�.�CFG7)��Ge�R� �w^�(�d�&��Ũ���]�@�E{��#\tV�?��9=>��0|�����|ue��}��a`����Ht���W�G�J^�q+����^<%�e]FɁ�p*�ܕ�v���v��z�ۃ��_�~Ex/�$Oe��/ħV�c�.���7�y�!����X��Q�2��;���B�^8�`��%(���~�Gt�;:�]���2l��U�3�z�3�'�˹�����yO��_~�7��N�|��w����ݔq9.�}�=~��~��G�	�q�J5F-+�&H�z�ʶ��xR��p�8M��z��$1'�^e���SL�GDx�+�l��	��ߤ�$��>M��B)�uyY<ᐥe�\#�6�:����g���2��Ee�M]3�ԓV�� �+|ԁ�~���4^�C��A·1X��>�ck������������8�nVi���O����Ę��kR������p!���',y����rn[�]:���"⻉32N$Є8�:��Pcc<�%M�>���D�r�Q+?�ې�C���g��u��}�3��c�{��u�U��fY�����v�
��T�����3�����0r����[�m��8U���/��K�W�>���Dihg�  K�I�M�(P�2]�y1R�`���8�%�[��� @�A7w���������T��o���[����k8��9A�{Ǻ ��6n�����I��{���
��Jt��-�E�w�e����L@�.�hD�M������>������.Q�
��Nv&OϽ;�|��9�
	�z!�C&ԩ.�����A���@�Zr����g|���|��GgG�j ��������9�N%�&a�(���"�{��h�%V&W�3�(�%Y��l�4VA�F��l|���JT2հ|��xL��R�#5�0�D��~���s�B�����F�Np>����0h;"��G��Y�{Q�+���ųb�5:!h
�)h���d$ƹ�o��pN�soTz��.�ܸ�r�S�����"{d!�A�k��{�lRG����U��?�o��{2,X5���CR�/���������G$C�Wb�߸���z���768e����	[���˗����w��wˑo<r��ض7wE{�)�Sב�:��%/_�nxf� � ��8���=GvASZN����
#����)LOMʘ����}�>��s�(ƇE�K�s���HC�_uC���+3~��ѣ���諧ދ~t�^@v���� �7���j9�l�`|ҷFF'�A=㒲�ss�`��`l�VY1�i��2��&�/t@ʌ>���H�-S�8��6�%���O:������ƙb�c`�(�g�y�þ��h4y�G���]8	�0�p��.���"u�I�Ĥ���q��U`�Iwl,���o��&Dv<����'~v��D� ��t]�s��zI0"c�ǥ���b��T1��N��g��qK8������EoR�vhH�zDڨ��$�;���?���Sv�u}^��յ3�K)�����	��Cv)3�I�w�J�O����Hp��:��O�˓�'�UZ�E�k܄+� ���^�MI��i�o�΀7ʈ�- 뇴�C��XmK฽�J��?�+��A6��y� w�8dp݇�)��8N�:a!j~�a
���;<	�0����7Dx��Ҭ�e�ʗ~>C��w�Ry�t�|Љ��v�������td�Y��� 7�R�>ř/e �(»��H�A��e `��A�a���)q��ĥ�U�5c��0D�R����CJ|�}_�`O#�h4��1�X|s(�*R�92�#��Px2��]|5B�T1��NE�8�>�z*�G5&}�����0~ކ $_xAֺѽ�je�
8���OE��x�� �́������^/``!:���(�]�^���?`9�O��Ztw`������ 
~&�.��sJ�3x|Tz��+�������qH���Ɍ.����h�D2��1NNX�|�8�������Gڧ�?l?��g������o�~%��ݐa;�		+���y�%
��v>~�n:����si��O��c�H)�a˵'�p�ׄ��$R#N�X����e��Ŋ=���O�E�}�i{��m���^����G���}�VWw}���g��藠�K(�ثIu�v���>��	�¥G��r�BO�Ȭ|11�x����x�B����לE�6��+ & )7�Τ�G��u�u �UD�[
�����Q�٘�2�)��uH��o��~u�2��(�� �x�-t�Tm���Q�1�N�/���wF�?�̊����]p#K��z�΅�O�K��x2� ʝ' 7��r��G�/~�C1n1l b9��)�!���Ǡ�^�y_eg��C�H�U�5��%��ܻ��TWx���D>	\:W��/A��F,oݼ��W�-���w�.��)�w�~W�#_�����43�ʭ����(OTN�eEҟcS�?d��/��arC��jr&6���h?�Qu����Ή�� 3G���A6��_�WZn�[�����&ap�� :}�B3����r�ru��$��
�Zл+!���g]ƹ���$K4�lJ��F�U��@�<��L�������u)L���'f%g%V/�ώ>@Ni�.#�t�_��'� %��{V�C�R ]3� �a{"���dO��B7�83���S~�z_���ۆ����ߟ�(f0��Li�E>��1D�H�rm��.�rf�a�Qd��c(@�ߔ?2d1p���-�/Ƈ���
@9Gi�Pb��V�ˠ�흁)�G~�S9�.Вwnm����s�"/��]:u	 א[��tF����=�����(N���K2�_��f��7�qO�h������?��>�����û����ާˑ`�̲*;11.`?&��6>�qyn�y��/�(�N�����_x�ږV��ށhb��(H�}iԲ���g�2
Ч��$F�L�p!�G�|N���~;9�~1�ĻWy��8d��������?|�VV��Sa�Yί^m�G_��^Q�����!,ˌ�	c�	U7��]����zH:}��ŘI�u�AZ�'=�>���>�G&5��*L9��G�L#�A���ώH��Ȯv��=�S4r�_Z��p,�t�r����n���(&��	(��^L�-�+�����W��'.�De�J��z���=k����L��|�{% �笫4C��1�Ԝ�Q
�r������?�9|�K������1��(}� ���l�!	�ˠ$��ȯ�g~�����d�{W����%]àg����F�Nx����#'˒�����ʭ���,�����N��rK[&<�C�B�D}H�tꈍ��)�*\���O�V�2/��� �1V�r���9v¢� )��C!����p0��WౢF' �q��s�u�
��%M�RF	@��Si�xpF#�ҹq8�]��F�7w�V��3�(މ�ӻ���\����\�v�/��]�;�璷��;#�'�J��Q*4�耳^�q�Q��8i�g]/��gȢl�*Y�7.ߋ���5�Y$���x0"��]��$UUm�.@���)h����=+h�bU2���#��Mu�VF%c�E/1.3N�?[��w���.@e��0)#�ݭb}�ɰx�&����V�m��/��5����q=zFQ<v�0�c��u�0r��� ���F�!�����>���Ah�Du��Ӈ|�靐�.��F������M��c�S����W�0=�Ku|9+�f�U(�^�D�g`o޺�-���2�=mkk�6D��+��d�kW�KV0����s����!�ű�{��S�?V.��oP�
*�
��F���/q�X>�&.-'�������pO��2�����������v����6
�
?}� ޞ�o=n��������A����	 �셁ţw��#hOZ��P'<��(�>��z�1�z}.th���NO|D�H��.Ǔ��b䡣J#<�(�Q���C�/�P.��۠|*[eR.O7�K�=�����3����N�����:�K���Hɖ�?�0�����R��p�����۲߳tsTDy@:�������e����ȥ��x�1�U��k�wi���|h6fƘ�(�T�����1����A��%˱�e��=\� G�o��g��oCA|�}�U>ԫ��:^��u#�=�(��qK^6"�!��.��$�ģJ
2\F������ۍ[��Hޜ�������2n��$�;��e�^��/��7��^��V�$�����ҏv��=1cB�4[dt�%e��A�`��� f
����>
Kgt�<ިk�l.����T�IP��T�f��b��t�Ώ٫����J�&�~'&�ȸ"f��Ǝp�L�p*��t�r�&;3F%�BB���,���~7h;"*�.�t�!�H�+�s)��\���%���W�r�S�x�*���Ya]#KՍ1�t$(i���AÀ�0F�Tt�̞�$�.���i$L�*��ڒ�Wnc�Gh�qLe�>�j���*�G���������z>0�<J?�5X���XE�S��|>�v�#2@�(���}{��*:���ʱb�Gc��nB���O�C���5�H����3�+>�E4�O�v��=V�����4�Bڴ'�(Zc��zD�!��Wa��䀤�I�ԙ��7���eCO<������XL0��%�8�py�H,h���G>��}��9y����ȸ@}��>�i�.��0�Ç�ۇ��KR�/Ͷɩ�$32����~[ZZ���տ�wmG��?Q>κ��ݸu�MN��[�ڋh��}>����/�W_����v�}�%���/�n�3t
t�l%>u�J�>�6B�$�ׅ*e����TM���Ѯy��3S�ڵ9���H3�I�n��=�LV�����r_l׮�hӳ���D����i��j4}<
�\�~p���i/R8�O�'2�y���&���=��/\OPD/�@S:�;��:ɋf������X��{V�9[����4���ك��$�+�-����Ç'Ԙ8�d�� ��O�Y�����J��vߨ�0*�N�}�#.��>D����Uա��9����<uq��� �Ť�VD9�G���@�����1�0.�ҥKD�O<��_��>�O�n}�!�m��~�%"G���<]�`p�^T�w4e؂�rC�uC� 8���,�g�ׁ;��8��Ψލ/����2�u��|�?�"|�Y��C�d'!_�����ԁ�F����!J�Ga�`�z2&9.�E�#I9���L��oձ}5k���v�䍶"��'���Uv���G��6�����#���^����e�ƞC���D?������*x��.ό��wo`��?ެojƸ�;�g��DD�bD�q������ND��{&�ҧ��� �����\���$ÃC�Qr�uccG$<o��TZfwf�K7��t�� �-��Fe%��T�p�qO CT
6���J@�ZH<?�%K�N��DQ�Ļv�]|�����h���b" ͤ	�v�����4
8�;|�E��#�`L�[�]��������qt�F�5q�E60��e�6ɚ�FK�%�ľN ��I�k^{���t�R$/v���θ����[���Nq�?V-��C�m|���&&.�iSS�o����<��{\G�/2Lh���Ȱ�q��F�`���.�Rܹ�"/�����n�^����7o0�&D//'�Ź3��-7T��E�Y��(�QE�1O�E���0,�6�.�����-��*㖶$Mb� l���ꈐ/��'O���ΡMrF_�����1�gw�.���c��ǿ�������I�Jr�p:p�>rj�c�T_��I�=˳��۫�GmZ/M�U���;�ν��k>�#�D������g������?�S۔�z��������w�V�vc�M�`��&�ţ~>���W�ړ'��P��H�U�৳6�h�����LE�W���Z��0/*�OS}�A9����'{\�N��GG{�c��ŨW[@Nȋ-�w�v9�U�.�����Ҥ���MvT�6�t���e��#�\<���w����w���8�P=�bu3�

��rx+��'0T�:�����HV��)�O��h��LL0U��?�g���?��:(Z@/�)ī��9��=��� ��;zt�_�a��G~�*ʥ� ��Um���Ɔ�(I);F�(a��tq�d�2��2��I��my�&���x��1�k@����Iׅ'_�eƻ�O#����2Ɖ2�t�^���|�B]p`����Xgܺ�)*Ӹ���L��e�u�yIm��h�JY�v��]Q�ޙ¤�s��A��+p���A7}+Ƭ:���)g�\>,89(l�a�ʈĮ�<��UƭK%c	)�׉k��$i	O=i�@~#�"��� ש��N�E�\�^�v���@O�U<2��˸�����p`��o����7ۇ��Ŕ�� ��`h�0f��AZ��<:���W���A9?e*1Q�;
�Wo���p�<<:W��8�R�R�j���s��쎊�&�>��h|��Ε���`:�'k�3nJL���A�䬙]�7AtҮ�T�!?q�ۡDU��᜝����͜��΄
��``Q'C��L"��wٺV���H\���f�n t�J��s9���>
u��U���a���E�%p�Țp�#�x&�F�<S�r/[	�u�eq#O�#V�"'�yS����&���/���8�_��Q�>��1�0T0
��k 3o�MO'�"��.����*J����Ld�bX��m��G�2o�s�.�JŅ̩�#/o��Y��Nyu�U�c�5�6N `_�B+`�ync�� z^�m��M-��?�(��������Ή��������'n�T�1�}YAU�F��G5Ng���#^v;���[��ׯ͵��)͉N9�Ab@�����8�`#A�B���;1��u�����75=�._���]WUƔp@{k�h�����|��������O4O�q���v���v��5�n�S�[2���O�nlm��Vk����pѡ���"��'��~���:���_��}�>�Cr�E*3����>�W��4��73�p{g�����L�HD���� �cVh�w_���*����WV�G�T��N����/ȸmm_�����ҽ�vK��iɱB��m�8�-���+j&|�˟�V2t�v��Њ��
��ip����tV���Ⱦ����֦�{�|llF���Ni{�拆�'�vA��)���uW8�Ԯ�%M�؋�񈶆�8�m\A�WZ��}����~E?m�{x��Uz���cj��`�C[���?�� ٱFtj�LQ^�ua�8����=�����ν�ha�a�{9���Uh�˘X�� �˂?�l ɩƆ��TF������^]�G?�)�d��Q��{L�|�m�Yn���:�*��g��ێ��y~<h���7����$���I��c���Ȕ2�NP,��K+Y��ŨU?MakU��*����Th�G�O4f�q+�S�t�ƥ'��&���/�p��^��a���(�ʧ_Bg���(���4*�/�b�
��Z�a��OF��PW�bCxJ�x�>���qC��D��q���h��\ϕ[�o�$�0"E���HSV0�(�z�N�+�*!��K[ҜF)��B&�'�����z\K��JkⱐAWa��GIp��5 �A�Wpd�zv���t����������E�S�#NHÏ�=�w@B޸#�P'��J�t8���+�%�ծt����<�,�s�U#n-���:�RК�*��w��p��[�T������b�_���h���d(�E��B@�u���3����ra�ڔ9�'�2�"<�P�P���F|�%�~z�ff.��w���;s���k>�����1YZ��(e(b`�n8���{�4X"[(�12�q,<�b�:B�A����ƭ��V�͋26���S����Wmkk��-��<�*#�Q��(��J{ �ܿ�fe��)!�0n�)㖶|AF�F_�51(��z�A+�dP�e�T�~9'�=�<"��;mmqi�={*��/}p��4nOx�È�IW T���P����f������>{(�n�+����)����v�T��*�	��t'�p��^t���R���䧦&|�W���#q�c�\ҕ�����B����i/�����e_�.zfm ���=�Q~ �|���{�����2�RA!E�ɤ�N��ؑx�T}�6�ׯ]^�=�	��	�3G���Ѐ�]��1e�6n�K�����0��mN�S�Y�'������wڂ&Qk�2v5q���O���F�h�0?=ْ���Lz�䓏>lׯ�Q���l��}������B��[�9�	l`P�i��Z�2F~oWO6��0�Q[`�Y��������/�툇ѱY����DT璁��DrA�''']GG;*�s��ە+�6�=�^!��� :�L����-܈V���� �(��*=%��uH��o���R�����6�v{2����ʽ0)\�k�T'��t��L��-WD���m�����
S?�x{��r����,+�p�B��T���.c��[7����N�� �ّ��ێ>�+����B�����g� ô�0@o]&/��H��݉:�����~�4/$zܥ�1�.�Qs��A��U���G���&\,�yB�~��&�M��a�hgj�6JӸE�~$|a�[��ҋJB��
-lCE˰���l˕B�oz�z��%�W�=����O���C�ޥ4n����כuud't�̨��FA&��^sH���q��Ji��=n(��R�a����eJL���[1�����O��p&�q��rR�Yt���-	�У� ~]D$>���@х2D���F>akc��W%�u��=��J��0b_��]�`�;f�.O|��*]�B�QFP�ѐ����U������/A���hV6V���2��/�(7�U)�$�Tc��k�ুK6��F��V��R\ȵ�"]Ȣd6�IcT6��;2XF�G�h�v�}�����3S2��G��0���N�:f,�'�Z瓶�"|{�h^L��D�E;T��ÿZ�����a{�b�}��|����-.�GB'f��x4��a/�{�����������;�ڕ���Y�X���
-��Ql!���t���r$���U�tّQ_{��8l/^����U���;?��)��(��+�;���]��*V�d,LO��������������wd N��qR�ϖՃt��4qO��E=���dܫ�j�H���1��e>�!�z�_�X?�i����j��-/^-��=n�D;u�� ��߱�8Ҥ۫��KU���ob����H{����ӟ|�߳�S>��'�4n�7���īh�5���Q�DJ�����"�Ղ��J��l���_k��e{�l^z�ܶ�%�	��R�P��3ؘg���[mw{IF�E�����_����ޝ��g¢����j�hr�c:�����N �/ނn�݉t�3��j����cee�=y������޼�PV�A,}�6�d�aTT�Q�U��������7��Lq��h�S�v$=�?�&�_�=�~:���;����W*�1�&�e��Q��%ۭ���b~��z��^��lj�xr�4lO���XC���1D�;��*��u:E��/W!"%|݇��a� c��|�I��8�r1�ꢐYO)7h ���.5�zEP�=.�+My!��LL�|�����8J��qQ��v��].iHхSrߚ0�I>�_���8dDoQ��y#�2n=�8߸%/Z�"���-_���K~Ҏ�%|t����@����o�F��-v_߸��ٸ5&�]
{�q��,��u0� #d��X<�Vn�O�����UudGj�n�BedZpF��J�Pl|��#Drx0K�c�",Q�-,��/��@��:�10nu/F0n;<�Y�A�� ��P�-a�$P |�iظ"���^�r�
�m	6����M+�?׸����7�=*C�2m���Խ/� �<��Q�y�sa���0j�RV��$Ь�a��)�������
����G���q��Z��z��3c<�ߘ��6n��1�S��rco�ф�-w�,C�\�����_����1a��>>l���ʕ����o���'�o�����[mB:�CL�C�g�K((R�od�^�o{�w�%K����IZ�a �2��񛶴I��׿~������a/�)��AzN:���mff�=|x����})��a�������wxf� .T,���%��5�,��)�l�)��{��$����~����h�k�����������7�̫�Q���i�%�i�<���x��p_�=T����������7?��{�]��=�Ôϣs.0��_�#��_7r\�~��׀g��C�D!�:~�sݗ/��?���2p���U�ۃ�j�h��o�-���EO������$D��f;�DkׯO��>}��O�뿑�A�~�R������ʎa���s�����0��v}���q�ӎ|n���#�&0d��Zm����~��o��ʶxd���[�_��J2�z�6����v�ʄ���o~���w�����;�v�G<�:�����W��*�I�"���)��*&12���	�g��Í�����Vx��&Ux���������vx������1Vo12�Wu��$�ѱת����'�������ܺ�f��h@��T�Ŧ���Ŋ<���:�&���5��qK^�藯D�;��}muc�=z�B��U{�������Ic�&"ݗ�$@������
�8�p	��p��-c@ω�����З��������]�lmtY�#W�D�q�\�ui��їb0a�b�O�GV·z��#v����s��B�;��>����U(�W���
��]X_��;��J ad��W�䝶ֻ�[�( >�+x����d�SqT�ԣm#�JWȂ&c�1^���'��Oj�* D��~�q�n��i�g{nܽ.��X}/��w&@޻�v
ȑ���Q*�Y��+�B�WN4կ�shQ3��צ�\_�gA�H	�k�'�jAW�	R��7䒄�&).�e:&�Ԏ��࿯z��0M�ʇW��ʝ
�9Ғ��^P��+C�+,
�3qp�V'x��`�8~�!��3*=�O�Sd���ݝ�6���^���l�����}y�:7>1��O|���~\��#�H����i{��(�B/�V:	�u.�]���ѐ䅱���cl����d��_8��7�1x|���M�����߇�Ȋ��?�N�a�0 *�UwV%��H����:B(����,٩6���6o����/^��oP���$�e�C��
��G��x��ٙ	���a�J� rL4���?��vɡ:౪��F'xN��Ca6�:���I�2tHE'� �0JR��8ؓ=��h%L�0(�v�mԥh��x��p��vI�N��S�!�pn{.% ��� �O��u���
��P�1ʙ�iW�O���.�[����W�D���5�I��&F��bt���1�S�Q�nF�&Y�c"�*;��3=.3���1��7�)�\u;!Z&1�u=����
6�P��	�*�~���.H�Fe�ζk�f��߈�7M�)G߱7^�qb������b�ݝ��hW�$����m>�,Y\���+����{ځi�vunZF~��M�~�pMp��d�q}��D�N�]�����v��t��p]i�.�g��&�IP�������S����>�}�N�F@��AZ �2�yq�t��=>)��)��}v��^�>q�W�^��'�
���Vu�1��"��,v�~�⃶�΅L�nt�.�A:';�����~�.���L�]�������WٖEɤ~WH�A�}8P��Ϻ�/,Ű|�'l�-�� b�-A��pN�\9E^DUZ�2��(8	1�.���帨,��'a@_�Hy������u]I�<�s\pU���ߠs�X�V*Q`�/;+fge�do{��Q�:Ew��ۨ����)���rH׿˽��>��4�$!�L0+�\��4t���mue�}��7���ʟ\]\��O[mgg׆���m�Ύ|�
�����������p������kۄ��Ξ�c厁B${�M	��/9����"S22��P��jc�Ϩ��ﴕՍ�.z��D�ʤ� ���=�}�{�ۢ�v�������ޖ�����B[X\lk���c_e�.�d��8��C�T��`1��A7?t��^uc��x��-�b��qii�ͿZl��Kmqa� X[�h|�ks۰�ے+�: �����遌z������ƺ��I� �����z�%{ak��?L��t~�ذ�'��������o�2�'''dȌ���ߍ�@������}诈4!:��H���R{b%��C���'2���1����6��2�/��xFFմ&V�'ե��+,����./��Xm_�J=�OA6�@\��Yh��;H��?�g�jWG����U�&qL��׵�T���;�tȋ�~�B�lM�D��6{�	�f�C�zb�F�]/LY-2�Y��U]��~�/��J דc2�y�,�-,�^Y'���^��&0��kN�`�c�	����x@�yz159�:PنI�0��e�j�T��Oq;QG�A��M�DP��2�w���C7}��Zˊ}��i��4�lr�v��1R{�I���S2�Sx��a؆q�_�b�,t�$����@���(��`�����9���I@�!z�҉��˸�P���b���Y�s��ގ������?�G#��������)��pS��tU9DyU�{u0VZ*9w"�aw��~e!g�C�C���$�7h8a��:D�P�/�����A_�#	��d���4,�W���v\�!/��'�}�;w�I��t֑Դ��-�X�������'4�B<�ׅ��,<=�S�x���@r�)��ʐ���3�v!�
�k���Ӌ���dX��w&�!��� �0l�v5�����h��KL�4Г#aCݣG��?��?ʸ���i��pX>g/���A��n(N[(8�p}�~�L���j�g_���`(	/{>�7�d�m��/e��Z��)ǈE�y���E>!���}��%��l����۞?_��;m��m$��É
G�,'��E+��_��!����A.pgg[�a����6/�vyeYi��Ĕ{Vj9�y_*'����exnJ��ƽ]�]�n�Ч����)N��i7o\m��]�zIr���f���ϯ�G_?iϞ=7-k�k2�7=�(�i�Ɇ�}�c�ٰŀ�G�ƭx��#�𬮮� ܐ�Ş�)�4H�s��k�������c�2Do�d���W�fb��#�6�ޖu"��h�q㲷`<��}C㔓VW����
�r�!��2`1|d��E1�ᬢb�ڨe5=�(��ߺ�5��X��G�ީh��X==���仴��^jҰ%���VH7]�ߕq�GA��kwn�h�o]���%e�/umoH���z�l������q��-cE����dɊ	���G�e�ǫ}�-�!ݬJf���#O�8=���c�2\9�cC�Q4�٨��yyn�ݾ}Ep�݆��i��<e9���	�d"� {�=r�A��%�uA��z"r>Є��W�x�E��(�0X���}�ΟA��T_��,1�`��}��Q7ԅ�����"����խӨ|���Q3�%So̧�s�&-���k��ׅq�%N�A�,������3�3���q���Cdt��%�U�;��u��_܇W�leU�*/�d&���~����}4��hx����@�͒�,���'��!<�*����:�7ǉ.��'\Uh\�&&���]���m+v�e�'��E\��]=ӌ<��̈́��ljϙ�r��B�d"�E0�����w:gI\�=���T�>q��-������!q�кl(��=iHƍ�2�9z�d�Y(�֔U?���t=|o!>��oC�3�g��U�N��[�ꀈ�WY�a����u:2����F������ໄ���I���p�p��)B�N��v��N�q�l��������+�$\��=aL��o�������-�/���=�OjМ`%���D&^}�U��o@��(��^>�	��a�\v�.��׃�n�>Ȩ?��CV�&�|b@m�3s�5��Q�/�e���+��� ��2а*�-Б�0���Q[R8b
�d]�^�z%�o^�жwo] �V:4�u�i�c9H"�_�ɛ�~a� i�p��8&���r�Z�����kM6���=��DA��`�:�Qw(�ma�tg��UB|�z9І��lnn���?K�K��.��*�6d�e]`�˸�/ć�ݧ�C��W|1�$~�'���X��qi��F+��H?{���P���mz���95�t�c(�G�,\p�����
��J�vd\b�"����'��+�L`��iE��c&X�L<\���ۈ�]&�.���S�V3m++�+�B���WKҙ͘tP�d {��v����5�z�`$^�۸L�Q�䉕wN̰���+�"?�G��W�[ �h���0)a���7�z�+���k��9"S��5G�.zI�`�3A�2��#��
�^I��.�Ɏx�)ʢ&��Ʀ&����]�B��A��=�'���A#�� �����u�2l���>��=x�P�
��{G 1%?+�� Y �=茜ro�^����@; '��v΁oq�U��,���p�G\qc��p�����5��������{~�'c��9.#M:ғ3t%��w�(+�\�C|=��k������Z��N2�N���;�e^���ş.�q��H�2J��!v�Q²��p��<�-�E%E~2��@_и`��D���gc�߇��A�Gザ@�F�� ���P����@k
�r��a����aR
��;���H��e�����0�".�ƣ�1�'}~���/]+;N�����w]W��U!����?�d|���?reNㇾ�s��P�B�d�q�+-���av}Q��@��9��˸.Kw�П�p�h~�RY|���X�bui{k�-Ȩ][Y�az�]��k�o^kwY��y�ݼv�]�<�Y�l�����(�m=Lϴ�3��ʥK�ڕ�vCi��~Zi�s�!+��|�e'V������*�y��8�J��GR��9{Pym�g}c[F��%v'6'�]��.]�ܦ�������q̵}΂��h���@�����͛�Y=fUw}}M��d��,OU'M���2��\�Q�>�Ad�jcz$��Q`y�Cw��,F����e�.Jn#���k���;�ޝ;��իmN򟙜l����!Ót	�����sYu�>Z�3�L��,/.�ھ��( ND�����ʈ��r��	� o��A<�/O��V�-�EFa�b���cՖ���H����p�����yW�*��)+���j ��>h|��F�D~�/���B�\�i�^.�ʷg��ڟ�G΋r��T� c
�[�°]�+֊g���Ĉ�K8�
9z����zԞ�x%><nL�MLO�H�j���I�9��{�)[�#yq�MS��2F'�GF��;�ON���T��#�#1�9��S-01b'�O��Q��c��t]:G��װ�����<!@f�����{&�q�%��/��^���?Yr	_<
��'!+k+��o�?~�u{�:�\e&,��F[�����AMAc����w�����*w�9^�B��/�#E�e2 ����@2(�:�7�x�F~���em����{ڕ2���3�#���G�)�F���'��O~����1�e(� �z����  ��IDATQ�[p=�� d���N!#��l�v&]�_��r�WN���N�]z蓳M����7�f�G�v��n���%d�49̉�K
��tA[\���r�w�YF�^��u��x֑��Z~)���#$h,�����Ht�9(Í ��HBM���girU�A��t	���a��p�\�E�+��Ñ�X����a�O�G�r�G:Mk�e���d颌��e��3��0D��.�,D��*7��t}+G�gB�+%qy�*��9��~�@��+�f�ُ4�!!���h�a�a��<`�8��ԃ�w8Ӛ��8��u��B�t1>�1N/�1B�N_jW���_��H��<uZ�xjd���ahT���H��'lT���a�^Kwr����1�
t[N�Ya�@+X��{�YMS�Jƃ�V�ا���̬6Q�r1N�ګ���lb�b�(�����7o�lss�݁z����iU�1lb�`u��tn�)uC�Z�"�FJu���I����+��l�ؔ���7.yC�5�We|_��iS�i�NSyK��*,�ƣh�$x��G%�7����>:���5��%��h�#�W:�+�19�A��]0 �U�TԣۍW��Ki����j8����w��Ki�����X�/�e���~^>��1?�:W��G����=��A�(��
�ŀ��S8@�]��ĦW�M_��h�U�^-��u��z#>����%O�0n��B�K0�:cH��:�,O;Fe0L��v��B�o�I�.ɱ�b\`�֙���
�Y[�)��O�� �~�(5yym^� @���S����J�JɈ\�k�F�J&��`�Ϫܥ�%Λ����s߉L �H܂2 /��r�;���DD�������r�@2.��i���7�?�K=�wa�Kv�� #$��c���kW�d��&�]�m���a�>�P���3�����N���W��}�7)�,�@�A��vJ[�Bg��{��+�������(��KZ0��y�\N��*��x�B�%�*�-����K�=��1@������w.t�_xF�eV<���_���TƨP]��r�����s��?����m.�����e�0G�.��$��:1L�0:iXEŀHx�{�*;0�8�N��8��g����L���ꮃPC����H� ��u�\p^Gx�ߏa=�9�K��Ϥ��2�0�n�7nɸ�&i\��#6�`u/V�x��pO��߮H^���hB��2/���M%ë	�����Ty�^{cנ�x��>�u�:IY#+?b�pŋ�:G?�P�3�:c�N��Oi��r���ܥv��m����_�ߢ�chF�Q��c�JY.�����+��b D�<��A��ңz�9��AF������?����>d�=��Nr�=�)++�4�2g����.���%�o��6V�_�xm���<��n�]�F�$���u�L}Qo�����⽦�	�gX��?=3�&���T�1��e�h����=>Fr��U��U����+�F��c�I��D ��#�:��� ����'/Q���Q�W�ߗ}��2�j���~b�G081��B�àNc��J �p^r����M�������Q�l]@�(3��x�xH@0�<�l�\G��G��]����ھg����IǉC�Ӣc����ū�br���ܶ��L�&<�b����_t��t1A�9 MR��P4�b�\�VT/��m8��e�V9E��[�'��h��O_C}t�>9@F�mt'Hz����w�ۄ%D]5�v�<g�����!���xl�tm3�G���,tN�[k��SD�H�U��-xz��?�%.�u�]�����.mp�¾����wя7Ո�9%K&"]V��JX�!��|��]��F-Hv8��������3���?ܝ��]άv����$o��U�N$�_^��a3�C3\]>a6p݉e�0�(�i#�0P�}u^��$@�)x�J��g��Ot�+@(��g��e��UNo%� �q�)������!4��i�����W1vwx��@6�b�o߯�	��z�7��� V9Y�3K2l�����21x�B�Wm15�!kA�pr� Ǡ�U�Uo���a��}�K����"����Nۆv��_��p���|m���ꬨd%�D����O�&��h���،x�	����$��&�Ǡ��_���w:�>���)F�X&{����^6���/4�7F�W1y�p _�~��ɴ`D��H���p���Wri7�iZ�E1L��D?=(JF>dK��9^�-䧞c"����O��݁^V��Z2�	@=%�G�ڸ�"7�TQ���Y���h�{��"Ь�|��⾄(�Ls�A�51����1�a�N�$�1b1R�K{�����7M=J��
?9�@��9���#�/�$T�ݴɝL1n1΃W_���6|z�B<��eD5C9�k%�	� Â�D�>4�w�� �S^����
�ӛ	M�XQgb����:I�	���`�:�.�
P�C����'8
�^tPza`��.�?���.I�CY6	^������Sy��Ҟe�����N"7�~�ώ�����|�8:���w9���\�s@�w!��tg��͇���3���H�}[���D�+�.r�o�I���V�}�J�o���C��_≕�h�(*�2͟'��v��㇋R�>�q�?n�˹���?�}}>�9��N ;1C��N? B�CrT����9`h��(5~ܨ| :/)E8�	�Eq���u'���Hׇ�m�^��:[�
B� ��dlt��*U<�4�c����̫+낍����V�W���R[^\lK�ŋV������0���sl�Mah��ecd�]�=�`�zg�zP!�"o5)Ǭ$*T����p���C�lI�Q*�f�����Gmw��WV���h��.�Q)'� ��8N&��ܴ1�=�Ցt�6�i�Uj����b�P���A�����[o�P]ז�"�\�Ȍ�|[����,>�5񰺲���K���mmmռ��U�:\�KP�^D�l[���	�_<R֭M�@-��쁞:�z%�۞��w��1Q�g�aE�/cFW�>!p��Ueo��4�ڑ񾻥I�&'{2����v���1�e�x�2)~�Zé��?+�Bza���.=�J�:e��S'����Y�1/9c�m�v���	\�*l{Su��g �pOz�'=ޑ��b���c���aP��mr����� S:���CV�u�?a�l�>�{����#�g���w����#��C���ɬ&����P�li"��.O�4Y�lS�lK�lj�c��5zB;O�̓���ẗ́��p$�E���v�J�a#�+��B_}-q�Ơ.W>m;簤��ku����gv��q�]��Ç��A�r1q�3 C�GnȦ��r�.C&��NEUP0�s�������F�t)i�3֗Ad�˹���et��;�=�)�nȩ�>z�[3&�	�Y�;�����rC�2� ���B�))���4v��t5�unp�>����BC�	���<����ȥ����ZZz�^��gڀ�ɢ�"ujC��40��L�Av��v�P'WNu朽N��rL7ƛ:��x!���"@AoU?���).~i^��O�6�m`�zL�*�BK�2��Vma0qN�_8�#�2`��8��sp+��N��Jh�� ��z�̒h��+��r��-N�B�K�e�
�%Ld����LW��͊�hK�0
�6��Z[��k#1E�K�
_��	��PQ��L�i��-,���|��x�^)�h|y�}�(�^���hK�Ѓq.�#vmͫ䝼;�����6�N��I���R[�_�$%�뭕[��>@�QC�*����fKg�eb��^1�����ڒ�a֜R�1��6��9|��޵�5׃'#K�6oX^�W�,*�rې����:'���9���) .�F�����i����"H�Ԥʄ�@Q�:��-(��E8�\�X�e���B���0}�&"[QBa�b�5F↌E�k�.���X��
��Or<���yd^[[��FBꟍ4]{�a0��?WH�,'?�a���8��ST�=�-��n��\�=z�K���yo{�F9+��!���#� �A�1��99T:rpmP��{ �S�k�괷�@�s�?�X��H��'<�q+�� �	�����3Mx�O{+��Aǀ�?ّ���C�WNe0Y����sU��F��&,~b"��hԦ���t�g]��
-�S/K�ay�.�]��o�tA���wT�Z�y�OG@��P��p����D*~ \p�;p�y�p���*}���q��u׻�7�?�\�ٜ�}h���%+���9�m���H��F�z�W(�.��@m�u�jO�������npT>h�wt� ��I�ަ(j��xʶa�a�?+#3K�3��rJ/��
+�~\�ǵX!/b�cU��U>6J[0h��I��y��� ���J-�.F�:���/eU���4رR�I���_����Q?��s�2����Yb��t]�|��z�$+u��qF� �+D2P96��V��Q����vt���P�U0X���+�}��Y{��?r�P�������:��U@�HgΠ2��8�j3Ǌs<�tR�!�awA2;�	Ϟ=mO�>mϟ?M/5�X�Q�##vW2�ۑa<�%��������|{��y{!X\XT��xD�#�cV�02�%��̓���ʨ�z�UN�6E��z�'���<�{&8�!�b�-���O�?~�������#�7�<~�u{�������c��Ӷ��B/��¼�v� �Ǘ��O��1�� �U]y{�zI@�0��I��|��E�<�d��o�^��|��b�s�ţG�D�c�So�����6�49��d�+ѱudS���X]�_o+�9�^v8�N���X[t0l��A��2�R� �����%DJn]��.��c&;c��`Gj[6`9F��;�5�X\T;	X\X𱁴�EM���ڊ`Iu�����i����@%O@X)��YC�(4�~�?i�k =��G���� `��mKNx���z�v��J�[ 6�,d��f'��^ڭ8uA[�Xy�0������:�ϳ.��D��C��T.R�_���<��h�Ј,hK��x��ϣ�\�e��,S���E����,diZ��/��\��|�du��}�uh���}?'����~y ��h*�|����x.6Z<��KCd^�U�.�Q�XM��@8���Bz�dqP�����W��D����Y_ux]��V����3��q $]��Owd��;\W0�g�E��Δǥ�Jڑ��!�H�*��ɏ�E�0�0ǃ/p����*]����AӘ=����R	���?#�:I$ ���I�;�F[�s���Nq��t]�ģT�8?����Q~p8(+ʧ�on�e{�<��䃹˗�����˾泪�f�f��:�=2����e��x���v�hp��g[�*>��AM�ߖ�qA�x@1'��>ӊ�0��"�[�ۼr����A���8.k��eQ�Z>:��d�N�L`�U��%~WdX̿x������R�x�bP`��FA|�N�����x�V]�7�X��?E��֫ggW&~<zf�ǂ�r�*�Gc�=��\�V}QjB��kCv�5����,��XYZ���)	��ah&}*�[$st�]TvzR�F�i,�4��|��.]�2C�a�_OەA�Ҟ�x}�����SMNe�j2��z��R��v��^n���n;9d!�D�-+^����cܲ��+�n�����г]�Fh��F T?��q5���{jPN�2��Fx�����Z�7Ol�8}s�4Okc��<*P��3�o�ޙL��	q��?q��O?�O}d�Au�Ne�l)�0�a"�:�hS�G�)��5�:f*���+o*}��ZV�Y!_��K;��<�'�(�$�U^&�^l<��W�ٖ!���51d���I�r��z���A��	�͸�2Q�.N��Q�3y�C�C�[[��C%[����H���~�>��m�
�Wy��e+>���Ǘ��gv��B.�D��O.�,�纞|{�m�w�M\��?��"s�.�{m�t��]$�+���
s萬�Z�~:�*=ؑ/�4�2������/(��Z�qu�-��z�����	�"*�
���s�q� �]�Y� ,�F�����TPǸ~�H
L��J"� �]�|�����e��%�\
T��f�)����q]x�w��Ky͛���fy��܃8�sM82�g� �f<;�j��,����>��٧�s��~���o��I��i��-��?�ĊQQā��+c��O ��z3Qu���0ظU�W�T?^S:��U2z]S&�+{�邎XaR��Qdt��O����p�7��	��6ᗍ�.�S�`�s_	;>=�q�ն�7m|�B��~�A����G?l��own�n�oݒ�ݿw�g�r>,{���ۣǏ�7O��P^�`�AP��J�1���/��?�����R�ԝ`T�o0N{	�1<�wK�c%�`��/�`�]�1�������>l����{�;�ڝ�7����h�/���͵I�G{mC�8[2xܺ��c|����2.��UV��\.<�����Ǫy?h���Ty�+^@�>b�p�k�wKva1�ƭc$H������#�;w����z֍k��ի��ܕv�7�9�JrD<6^[Y7�|�/-!g�qLe���
��K ��k�A[�Z��H]��0��X}'�9��;'i��&
;�y�|�#�6d�>j����[���˝��iR0��vYחg��M�I����X�-�"2	`��[���-1�l�H� ���x�'9�&�>�0�7^��6�A�`��z�"|� |�'�g2��*����M��S#���K�ֽ���������n�[w��+�fە����m�U�j~�����m�ΰ�}�L6m\���bh��j!�nG^��Vx�T�rW=�sL�D�/� �̾������vE��*,��^YYP�]�1>{i�����4�Y�gDs��#\Ҥ��8Rݭi���������Ɇt��6��0��XO�{'��{;��vfp_%P�PG��.�d=��}�� �\�~��41ʙ��s�>�q�Oś>�����TF?r9Q��>�^�t���?&��&�f��A��E���K9K�?�	3m���@�R|�Yo�?p���mS���3��%a�Sŀ�Y ��C�q�qL��+�h��ٕ$ �_�Խd����H�`W����t�/pH�,�ē���h?����`�_<���� �E���dT n�U_0�$���M>X�-~~��K�QV��đ+�y�����H�����7��2�^d�M������]��!�Oc8�Te�td�2�#c�����]�H���!��H����9��}�_&~�9��׃{�9��tY�Deqٗ$J�S&�!�uiHa��ȯ�BG�Y=Fn��b;�����89�:�!W�iK�2g\���H��/��{ȃA���xĪ��2�,��=os�������C�ڲb�S ߩ��*�Gy��ֆ�ϟVl�2P�I���>�j�6&h~r��b2VJx���S�����Ƽ ��D'G,1�p>��}UtWXm�����e����r�>e��pѺ��Q[��I�BWݲ��J��'H�3�>lD�x�)F��տl���W����g�eU�k�Y��ڵk��MI����5݋�\M��k2no\U�|>������K~���t,�	b�|X�w��;Qk�=���y��\�wq�.%U�%�n���&Tl��4x�y���3��7��x�&�]�Xȕ�0����w,/^��� ʃ$��Q���>r��u�o�

M���`��EFL��,�-7{*��p���W�fd��]�ܮݼҮ�P�\W��A{��t�ton�]��:�)l���8&5���������a���HA�~YQ��J��:�C:�3
#�C~<��d��=�[�L�������=�lj��Lt���v���v���v���ʕ���%?5�8@N����D���]Bx����>�ˡ�*pKWx����:K?^�C�B>�r��_oGP^�bY��BcE��.T�9Jz"�i;�e��x����k���At&ÕoG����.�&9����~�u��~!Oc � o/?�E?:H��:S����W�J�:'u ,�ǱN�	�B�IA���q��ҏ��Ɛyax}�3?�%��[B7D��48+~�QCi�꾃ԉ!�8��*+4?��?��.cϝ��K��J� � �q�Ho�/s� �"\���uxh˙�
�U��PY�	ǵ�"q\C?��q? W�5%_]��{���|Հip�	$>�R�
wY�ͷ;hC�=��q+`P�d����	��Y��f�`��x�R�۵��T���߀�L�6?RS��I�����"��[er�h�0 �m�����6�٪�.٘��4+�/���	V���#�}����d^FaU.>~�j~�=񲭬�۸Ş�')w����;����8�J�J��"¶Vp�s����{;�3�B����=?>��,��hQ�J>�Ni�(��G��T�KV�&��_����S0��Oe_�(��E4�7e������W��ȅ��kAu*T���i�ۥ��7���,�������2*�j|؁Ig��e����]��a�Wp��U�]�W���'U,�c�0�:��B�?�-�-/Hq4+��a�Vx���]O��@��)�?	+�bR%v�4�Ub��O��_��5_��vNw���Ӏ�{�~{O���ww��OT8cͥ��� �΃�d-��Bt[�"�+��t-9
/���'�Bg�;ձ&|^���)��iQoT>z0;�ɠ����9��mrZ:5�׾8�y�M�~V�/����G���X>8�J��۪�ė�x�v ��z��=�^�U�bkP�P��UH�4h0���R�^|�F��������g��5���I�%M�nߺ!��n�S'����N�<��s7�M*tM4��8��>��D�qa��<�'h�E�I���5��9�C�ZW^�.���X�CUW��|��|�lo|�� �����d�7h; /4�]�2���K��`��TX�_�������[\����+>��HF_?���\�ͯ�髻�0ܙ�.�W��*�ʗ����b��HP�0�w}S�}���u�=s�.����B��sOM���m�%�UB/���}^������e��-6�+�( ���:�tq�S`����L�,=g�;i+q|�C#h�n�wtq�.�4@/�� �v�(��UJnWbmc�cM�� z�+�m�&b��>}���4p�!%t�`��]��=�{�2�x}|rA ÊGbJ cdљ�yQ�9�?���CQ΃�i����T�@�>P�Ύ�8.���o��u"���A.�ޖ�`�y�Fn%'��g,ȐG�����{V��<pA�q�iz}�i�#kN��8��`�8����?��5����M#��#d�C�]�d�ѣA�A��p�5h�r?�]+��9�f�k���O��Uj�z`0]��ʊ9+�S|�����/A
0l8c4Vԧ��X�3&C�_���pC@�����K�
7��E����Sg�"�缢ˆ�e(<ɟuU���V}c�Q;#���-�p�'V��q���p�	O���Y�U�Ӗ-3�����Ӏ䅵>��&a��t��a��4w�1`�Zi�J�}�IOΩt�9�	�Q�RƦ-U�k�	����)���D�ޣ�q3��(�$yr�ƹ'��,���
���	��2X��`����"�.%�v$|���	!.�"����.�6�o���� 6VlY��ڮ2���y��@�~�{�9dI'��e�!*4t[q��@7y��r�{t��$�:qݫ�\�L�2�EY�䑐�3"���c2ܭ���>*�^����}�_�С�+ׅ���&K�g"ȅ��}�s��
W_}0�~zgP\/�w����δ�aG�<��8�W���GH�����g��#���VX��w1_){9β�==�2gRaR��m`@*�!����O:*o�lYDU~�I�����t�g��9q�6D��4��i��/?d�_�@��>T\@���#P�ȕzG�8`E�AKNq$wN�c�5��?��O']+�68<P������=~�to>4(�gcB�a�Y�2�7�i`�-Bƿ��y�]рue��1�[2y\���L����(�7/��2G3a��Wg>Y˪M����9y�y�Z��j��*��#|�@�?�`�d�f?G>mnp�Ҟ�d��1���c������>H��ZXxeX\�,�s���v:{Z9��2���I�K^�����%�0�0�x1�,cѨ�9���FB�������aQW�Rc�.0T�ԈqV�ehO��*V��͊rNd�*^:L�����t~I81j�7*�� t�鰣�{��0���P+h�q�$�u4�Izd��?*�#�U:��pz�굌��Ӓ��abb���Nz�\-�DbdP�}�Ԇ�da���}���#g�B���t�H��؉�7jS�3�����ҍ�+~�ϜD�wԣjg���$ �!�
0	�i ��Ư��32
g4i!�G�ْ�9��mWr�~��r�3:C�9.�ഫ���#�^E��/��
(ȯe)����}MLU6/��o|=�'| ��}�L*b�~�Ǟ}�L�j����J�Ԥ&ǪǠ]} z&y1٠c�T}Zo�?WV�dt.�J���t�/cv��]MF������e	Tx�״��H�I6n黳���[���~*��>��a�F��[�t�و�m�a�1(��㹑���B�Hu���y(?��BкDxOC?B�v��+^���.� 컜����H]�`ȝ�r�z�u�qh�_�A۹��2�	���g���0.J��AD$�uw�y�������gs=Y����3�Y�/>�:���]e8A�yx �N�+�i���9����j�Gr:3��rN���^^������+��i=87��@zp����m_��&+�����V��t���oC�t<J��`�e/#''`���r�7�e�z���ZVCYͭO�b�I���vxp"#�m���\�h��Y�1H*�>`\*qX2����Fnl3���R�km��v�g������� +����|E�[�/�qL��x�6��Wz�G�Q�uD����Y�����^���i;�[�?�6�~f�$V^�6���ɘ>�GmkK|	�ֶ��N�3�ұ�jc��WE�;z�A�>UVȑ7���ˑT|��r8�-�{��<V���O�ή��c����6:�7��E&�Z���f����'�~8t����[T���n����Z�s<�����A�,�B����L�� t��:����1�54��������x=�|�sj��$��b����vn��f�nT�1�LJ0�1,����nL c��&Bjo^�G7u��K�\������|�#����J��=��a�T��� �'�;����[AҸ��[n��/��	gS�o$�d��mJ�7w%_��z��)�/}����+ejo�Ig��'8���&�L� ��.㖾��=�=��UF蟏$t�Ha�(���{Q?��
D���o�֦��4�K� E��|��#��J�r�Ieت=�ҔOV�<\��LO����#u�@t�y��{��,�Ÿ���u]��'�� �(�
����(��t�,up�/֏�+ ׯ����r�E�Ÿ�׊�K:z�����h��D
�E��D��z���&�
aE?ѡ�*���{�U
�J�������;�ħ2����X~����ѱ k5؊W=pDwO����<B���Q��$�Ew���Ġ:(#�̲��t���q�Ϗ
�.��V/����r�M�5�bTm�HXZ�hϞ��o����l�g϶�������+�#F��\;2\Y����Wۊ�\��qN)�X)ep���h�G���qf���f{�bA�>k�Ó���g*wY�Ldd�UG5����S����^�\hO�η�O�ڳ���m;p)���a�As��p� �㧎�a Q7t��1nOY���T��d2�9aEe�|�Ҟ>]��VګW��60ٻI��2�) �D�>�Huz�Xh�"I�F��Wk���˫�=#k��<!d<����=��D��+|���W��/{�H��d�������s�)�����#ɐ��2�B�0jc��=У�xJ�vN�����hvd�S��Ҿ��P��㶤2���m�Kެ��2�p�rL�m���-� MN�K�A��c�����sl'�3��I4E�̊kL ,���(�r�8��������wF�`���L��	�:"�4�鴭��ŕMet�Q����I�2��;����]?��'ɓ���:dE_��5�$����&%L��������gk֗�������c��)Y���?���0d�`ʨ�>{_�侾uҖ�O�s����f[҄s}k[���d\z�J8��ĭ�����1�γ]lKy�-G~q���ʊ��{Чffd�N��Q�[[2�7N2���<݉��$s�p"6�i+�FN����&Oj0nI���O��Y��d`��>�Q��{E������N/]���@�\t�!�{�1�}pV��W���"*��U�Y.�.��΋,�@�<o%�#AT�R#]����+>�x����,�+} ,'#�s�Ǻ��#]��2���F>�����9��vz]� ��ʙ!
l`0��+��D\����d��0������\�Jk+�3K-7P`A�q�2`���"�Z��>*��@�x�
�AU���ce*0��!I��e5�D΁�T&<�Y�s�9ȭ��]�u+�g!���D���f�����4����d��U��/���(q���ˌ$%�z�D\���]D�E�o�A[�'��8�F������������Y+L* u� ��ᱰ�^<���Dlg���69�>T
�������~��A8W�U�^�b���ƀb��U�M>3�{$�
�����km~�3\5h�b�ʠ�eÑF�Y4� ǽY����m�Y�!��dm�>m��#m�2�7L��	ѥ|<����%U�|�Jt#V��{K����n���� ��elR�i��ܓ�������U�c繺U���\$P�d���+�I��	��Һ�w�̵��M��c��b��k�g��t~��#f��I9��>AD`��n�췕��6/Zwdh�*|t\��/7em+k�����R�,1a�DC�Թ$��ӂ�?|��aǥxw,�>BMF�����6��������sI��%�7�eo�9^�❷��c���"���`�+cuscxC��jS���/#�X�s�gJ�}-݆OMP4)���u���?� �]�n�?��X�����Q�cB���p=>/\q�+���e�EO�)��i S}���-n72.0HYU%0�bI��L�%�2��04%�#M��8{Z�M�^�\����&A�B��b����$[B$�{}���jo��Qϟ�҄�p@#�R�3�m��h���.xI�3�Vmc��"}����/^�w�����v(�GF����4`�\����h���$&�Q�����F��L��̻v��E;R�p�y-@y��}�k� )���=�\|���J�]��n��x(��w$���\gO� "�	��+���GX�W�3����-)�����~��P�С��9&�w9�)�G����*���c�v�I��x4�$#�
����?�b�~E}hN����f�B6�����m;
 +��7���*ot���u�E�Pe�Oݩ�99rx��%���q�Y�U�
��z�q���5`� X�T߸%��~��NE�%���#b|M��E8�(�]�a��3D�;�֍Y�i�!�J�����E��c�Q����h"%q�Y�I ?�*n���e*+�'�;P���Y?^����[��!�*�qܡp��e�����P ��&=�EeL:��|�׸�a]z�����CS̪��HT�}�:��vb�{O�~p���������T��+�<��8�rwǫ���9"OO�Ȩ�a���Xm��	Z�{��AVkxD�cM�ul+2\1h�d4�o��;�eD�0�kF�w��ߧ�>����U����xVz�d\b��x��gi�u���CQe�N�k�#*C��%^l� (�p������5�c��H[�5dB#�&��=�k_��q��+2�9�}�k�%>� BEo�ag0ypf.ꈺ�	*��0��"+�K2��_-�L�Z���C����L���1ڼ�#�u���z�z,��q[������%���@���<^_Y�l�_,�g�ګ���ϯ�J��^���/&��_�PK�ȶzG%�>Ou0!ِ��z{�r�_c5���Y��c3S�����x���ɮ��e���{��x�?&r.J4YR�c,�>V7�ږx&#}Su8?/#T|>1/���+��ıc>6�z3Ak��v�a������Ճ�%�<�_�2���M?��nf��8�p�ɠ����7���_�1��3��� �����ǇO�g6�e�b$b�b�Ƥ��DKv�l��:���G��h��2/j������Т�����mhQ��8=�)��q�Zm�"c�du"D7/b����' �e�{�Fߢ�^�\4d�����jr����������0�B����vtk'�����R��Q���3j$�z��@�fa��Z�O�1r�B���	��Ba��^Y2M�/�o7�Y�:�8�	܎2�i�N�-|�_��cp1&��6��_ܯ�}�{�s��s?V�#_2�u� Wʀ����VGq��q/h�O���r�~Ӹ��	�{;�!�K�,�[LS�`�~0ޒ?�j�^���2�f\ s�S6V7�2I�� >4�xubz�[����v�]�ds�ӿ��[:>2��,0a6�3caD�`���YH�q����}�r!l<��:��@oZ�o���t�I�Qy����G8\y����?�%m��`�Ҙ�N
5N~�lx'���	w�/�v����> ��=?�E&e�;,�$C��°U��C��gd���"�]X���R���`���F��$����*��'��I���D��)ՏuJ���I���l�Z�PG�BA8V�yԸ�g[�ٖa˃��_ø��'cEm��j�cg«��!w��"T{9Ɖ���{ �<v�8\��o;{<.?���c�MV��-��`�����.�A7�,_Ԇ�'P&�M�n=�/�d�52�#�>2"#�U�K���bM�K3�QϾِ�WO�ᇑ/�a��P���o��V�0�0
 Vv�1yI�f���iCݪ��ƺe3�We�����6��D���|�=��GT�Od45�f�^p�:���PJ6�POÔ=��^�������{.ً��cQ����jGu#~�:���w�'
��.���p�v��O��:I����k�Є�U�|��-{��|�݂�+s���IM�؃+ƕ����pbo+����6���E;+��C<RW��W+׬�b�#�-�͞�˾V��`��a�;�[&���DJ��j'����U�Lh���%F�-�	�w��>5��7+��Uۨ��Z��0�7&�Ú�kMx���&\L�`82�:P8�o�[����cL�/��fy*�&�0ni�8�̓ɕ?3-�Cyz��8�L�c����W��M=��(V���NV�1n��d@/o�ɠ�����Ǧ�D�y�[Sh�ٯQᦞ~F(�8t=�� ���Ҙ W�%[�	 ʳ�R��8Cn����Bx��D���������E���.�~����[��K����(�?ӯ(de��!����s`s~�� ��K���#o{~ݼ�)���_�>����\nPS+�N��=��xL���!�Y��|����;P���4�'�PR��;d��@xx�T6V��K�7�AV;��mN��k��i)������q�nI����	� 0�A
2�J�̘
c�׼dvp��ڝ��# gW���Rt�ۅ8��Ё�ڒBPХ �H�Ļ��k���/\�H#N��'3n˗C��?p������Hp\��L��t�R�\�R�QO�s� }9*��Cu��u���/��_�{�Vb����,E�}�.|#�J�@�	"N�|�&����"�0Ҁ���ƭ�FI���x"�On2����(\|P��1딌��0e`ty��>)e����8�h_81l�4����(8 ��'É�:7������~K�`Jՠ_�*yl��t�:��i���쉀�]�	�33�mvv��,g�N�Rƌ��R��dz	Sl�`��M�܊n�	l�a{�1h��}���$�����=�.�
Q���"�W���������+�(���*���}s�/����>�B��L�*��/W��W������V�{�1t1l�B���yJ>�M��	�C�cv +�A�����O*�]W�Z�2l�n�xlGF��e��$9�3&����v�r<�W��R����z���3j�#aH�\XZ��Ɏ�%�y����}����1ڰ5?�"�m���Iה�F�>�@�ξfVYwe��$��s[0	��S<��ׄdʏ�/j�]L^�[ʡ�G*������I������'����Y��c�x�-������	��1�m��ؗ�1��#�2�1�1V�������"٥io��g��Ut�\���	{k���+��8���64�q���a�-=`b���#_��=�7�(�ap*<��D�u<_x�ѮD��%�P. @翯Wu��Sg��.��4pRvJ�6T�N����{�),�.�Sf��H����.W�w��V�sQ�6(�,@W�� �Bi��;B�x�
���#/c�IF��e��w9�(�֘���ƭR����P��,~��i�T,u�Bt~J+�l_	_G�/�'@N��xݖ�'} ���zT 	��/\�k~��'�e�q{��������|G
NH�t���h�a���e$@�|�p�����\/��q��/gZ��A���,���y��8�z��ay"��]?�<��
�C"�z��r�fw�cg���%KA4�j�� ������:i��4f�^�;c���Qn:_ihL4^B��&:D�\E���uN���#�x�A�
�ٲ@i����Pea��[�t`ʱb�ٲk^%3NJ�bq��(#rp	0sp��s;E��kR
��B{�sbU>2T Ձ��9��LY��I6�ԥ� G�$��&�a��^�:���;�c�d��X�q�ct(V#Г(F=�Ȉ�[�M��Fd���]��1uAy�X	Uݒ��}��T�\V9�h`��b�D�$��vD�E���B��LnR�؆�#g^��9V���7i�U�G_�&@� ����9J���N:�^K¹�n��	:��}��ꏭ_���z�6��t-����=0'qg8.LdIN�e�b��t��*���\�&@L�;�ckF���cv�|�'|r����bą'�\�E��a�#|����-ANr��ZӎO
������$Om��|n�4N0�$�h�Q/��d��,�Ř��c�2dEa|яm=L:&E?\��z2 c�m7�L��M:�
������/�Q#��J=y�pY��'>�B�s
��2Y�}HGfdŶ]�IҮܾ������[}���g�pF.`W~���x�sx����'(<��y�}(�k�}��`�b��r���;_i��/�A��=����K!^���P28{/�!җ�����(��΃tu�>��Ut�5П�h�e�`�.!80 e6�>�(~P�Wsh�OG׃��r�WUk��(J��t	���׸��Y7��㺼��l�}}p*��_�;���0`xӸ5�Hࢥ��e�h�d �b����.:�x�(\�!
�o#��K��^Y�q,�i�Ǒ�cmfV��S6:��RV�a����B׸�x>y�?���@33�TƬW|�\�ql���L'8���!��y)�`t�a:JB�'���<C���B>6<���`Ȇ�2F9����q�>��(��o���l���_~x���T�Ȅ�Ag��d��6{\�F���YɈ�F6p������5�� ����1 �N�>�11�L��k�Aަr�M�����r�~*��<:{�1F��~)M�PG�SF�j�:tSm!�������w}����? ˲�6����2}D?�+~n��(:�"As@߀�����hR��N�ġ'6�E�N1�?!v��W;��h�>S?�ol�UO�+� +=���1��1Ջۈ��1Y7J��W�3� �2��z�8���G�E;�="������F�},㜭1��S��r���C]�5?�c�%�vj���c#e��C�!;&���sʃ'n�I=�N�QK=$;^uG���	�w]�$v����DN�J�f�%t��	�T A9��I�bE��L��b� ��w� �rj����2��r΀x���K�ڒd��X���6ae��ԙ�(����C��w:Ҿ�/���B�]�����?�{N�Y=���1繡�J�iM�����h�4��`����P��c�ݑ6.�������:*�/���;/쇺w�����̆@rU��nv�w�~���Sxv��х��ŗ��׼��D�Z���)F�H>����9ڨN����! �sr��E�L�wtb���/Vc�'q�h�ȔU��Ł�H��T�1r�a��#'� X21���SF����J�&>�d�`Q������((Ð���?��Y��+Y{bL9���.��^e�q��)���Z`��u�\���I[я��d�A�}�@ܢ������aV�S>�m ���c� ʮ�PY��	��yɣH/��+�O�!/Z�� �<���p�L��w�E|��#y�2���l��\����O�[C���'N���!R���eiq��F0�';ƞ�1XO���޸&]��_�t�K^�o��.��<����!�>�OO�TG�������i
�8�e�E��w��e�Ӡw�E&��9��ڲ�#{����t	:��R�L��>���ݦ!��{eD�A=%�"<�/rb�N?^x"O��B���Έ��o=IJ�6��hML�9�}����\�].ˍv0�,��\�lP�sʈ$Q�n¸�6����tNG���8S�E[�]�F���L������y�S\�b��ƒ<E?M�����JnF��9.��ݙ<��"�]��3y�"H��\��]�	�9�K#%V�ޏr��-��%�%�=�]&�\�V��G�s�~2�:�C#�����P�������9A����:�����8x�!�SR;.�|��S9��mW��u��[������}���AG�x�ܙR���.z���:�r�Ý>'8�|wJP.��еz'�XE$.Q�|��ȖS|��){[���W���Zx|�<Ɯ��>0�c������ȃs��C��V$�6ԁ�H�E���k�!����A<rA��C�J�������N�-�_���Q�B6>���J���9i|TS>^eϰW����~��X?
t��h7v\�b^��6ք��0J� a�+���j�	]�/�U��2@�H�+nYi���B.H]�!b0�A�\pR�M0���&u
 _&�YGE�?,��y�g�
���%m������GpS�xG ʨ2ŝ�4a����G�%\\[F�G�����¨����҂��%m��J���J�0
���P�5qC�gn�XЅ��D%W�1n����ؒ�������%&��®t��.Ǥ�g�Jg���j����	N�����������X/�����K�w�Qw�+4�2t����ݶ��do/�XU��a_�>��(]�lB�����h���FB#�0��=t�u Z�M�e�-0�ӑ�������	e�l�g�
�������.��'8�y� �z�I�)[O(��dt.�r���!W���VY��^�Xzi�`G�gA��?ǙȬ�*C�����<�̂y�&���&�]?T@�~�b�VxhY���B�� 2�6��^I<�7�A a�V�/�����@C���d#�J�7s�֕���^��S�ιK�{?���!��G�c\�s�~�(��/�����tu��<���J.������VGu,@��3�q�����
�ԯ�v��\�OpQ����� �{6:�3@�(0�:~Vxs�0d�]��OMy��0	*�c���<RE�i����S��X֫X�G:�v��Y�t^J��`cX׆_�X:��@'��\�"��������"��+�i0��\t^u�2R��V>!H���AY�^�:�;��Q�n�+8N8:}4m�#:k�NT�΅�õ�ނ��Ε��s�I�1Րc}�X,O.�s2o���@��ϧCP��W��Uz�i&;Z���U $�s��ƙ�������Й��Q=W��"ʴ^a��Ot*tKXL>u��& o*���<�"F,�����3�¯��w��3dv�H�G�q:*��"ƨ�>܊f�����`�W�y���zu㗙Ƀ��O��b F;�~��ʑ�@I��`�ah��Q�����O$[�� �a�Z�-� cp*L|�	��4�p�JG/`p��@-\ ��+�E����~�}�d�{�+A�q�� (�C��!�"��(�y�İ�Ͱs�/y���.�^2��̷þ��q
� p�ύ������'>U���t�s�,�6��A�iJ�|���qN;��ޕ[P�_�]&@����;�D�1,�Ե�"	~/���o���g��.�9yqCu�m�O�:ȸԁ�/ ��y�9..�u)�r9�܏��T�y_��>��!�i`���Y8$!���8%Yt�Q#1TCQ:�L�k�B4���%�՝�=� Qfu
�;�һס#!LL*��*��х��g�K��O�j�@�A8ܻd::>�5(ĐI̿~�'�2dä1�,bH�������Kc(�%�"�t	�i΁�+�8�����:ʷS��Oe@@�B0����E��Ǖ�4��X�=$)��F-{�x(�#wJMܱ�N,F�db��D�q�J��	��X]�P&ر3,g�H%���D��%Ƨ���̧�]W��'����v�
Y/�@x�U�0Lx����j �zŪ��8:��1��w �˂�hF�A��aQ/p�αJ�2E�����S8<������U]�*ĬA'*�U^i����ݬ��ڔ��W�j�N�2ؓ�~UV�b��@���~��BD�|���+�'�#�IM�ɋO���c�� z�����W��)?UR��[bV�S�G��8��rSq6��7ݘ�r�В`i�\D>ieQ�$�Z�G'Կ����
�:A�'x�R��'�H�����f�/oI�]�������5Q�����C���>/�0ny��S �Bg:f�v;+�B!i��I�W�D:/d�� �8?9�!�Z|�}��L���
'+��ц�
��%��D0��T��آ�������.�L���#�t�~�9�8��Qx*�5G�q*�HzB8mH{�B��[\�]8�v�ۗ�L4c�yɧB|���+�'I:����cq({���~S�c�10���'P��/ �p�=�$k��6#3VCh�����K�r��VX���I ����.�I�����#z�K�ѷ�-�l�#�d�����UYf�(��6��L�U���%�V�G��t�S�;p29�	���	�0g<)�G� ������?�/\�9�A"�I�^:;�K�Я�%�%�NUǝN ��~)c����W-0�� !�.wN�Ut2 ����B�Jc8�!Ã	��殺�B�t��#)i
O�����r��*���'U1r�@Q�{倣~YaFY�D(�������lx=�[#���Z��' i��'��r����{JHx$�4*�<�i
4��E�s]��]�4H��׏�ˁ�� �H"n���V��Ye*O\�*�%�{�!L�1o�I��AR)/9�
��\(�vT��]��?$���TF����2�l ��P�Ɓ4|\V[xA&�o�1 Y@�P(��YN��D�2��I�w�G�b����D�q��O٣�=>���a���"& ,Vxe|(��2�&8Svz�MNŋ[��te�
z˨L�̌eϯ�������\AT�+�U$t\ :�k]&ꓚ�&:/�)҆`|�U��lh2�dD�/�%�n���3^��A	U`Z�	������sig�>Y��ě�+OĭW�
�L�d �����C�0^ѥz�}"9y%�3��ܲ(��'+�!^nb2�.e�1q#�S|�'�"��;F���7<`)�l�L̗���C:b\y���0�B׭_@�a�ԣ�J<Qo��O0�Lm̈>=��sl�P����hڒN�#dP�+>�k�y��2�@��J��7�3ȓфA�'-	�.[���S�'JK�8��������������f�� ъaQJ�2΀�+΅'@� ڜʰQHm�[�W"/2���0�e����������L�-N��Y�B�6�?(D�!(����{��	�2�d�[n �C/(�$�V�{���!w�+g�����ޟ�Z�%i���<?�g3�"�cȩ2�"�Y�U�I�D�����rA����&@��E�t�HP]9��>���<=���>9zT������{DV��=�9r�L�G���#�S?m]z��2�@�e��c=Dn�I��ģ��ʂ*~	|G�G�8De@�D�H��XO`�Q
/64�f�˨�`��r�?ƍp�8�ҡ�ϜPV��$E[��[��H0c������9N ��?���3a�^6"�*��w)[ਓ��n��E���왈=y��0�pAit��+?�F����NGF�q�V%� ^t|�D����Z^�J�F0�M��y���ҋU�y��%������)Z-�{y�<��Gvm�=۔1�XF���S���M�����y�����Ñ#��/jx�1XT���: ���&H��]a@N�lR��$˘�g3C���n�~���;6>z�F.��kQ�c���2*�����a�������[=u\|�"~����"�ꑿ��� ��v�_-Ee~&��(aA���{�;>7��'���6���nW�A���1l�Jg���Cn����]x���c��;Y��x":�k�N2��i��0z)�!R��ۓ�$>rK��բ=a�sG�E?K�t�>D_���qC 2�ya?�v�<�����c���~�����ݺ 9x�7|�ŀ�\�Jec�R.m;�ѿYB^w2�@����� �σ�Q���!/m��܎�!;����F�� 0F�C���#Q��z���Mc:�Q����S����0�	S'����!7cy1f�`�j|�_c�p���<��?=�$c��.�p�/q44}.���1���㉋^ڃ��b��{�С�:�HF���S�:�F�@���w���ecܝD�t�������`��T�����q�f�g���^Ǹ�ڸODw5T��=n�Ђ�����@�Vl��\���_Pzz���X��Qp�Y��mlJQV�r��e�A�Ot1Gd�6"��Q�B��$:�����4�cP�o��SZGA# �bg���'u��o�E���qXz��b��
�̛I->��t Ӓ��v ��T�R�%D��G�Fr��ճ��0t#~�8���f��G+�	��YRV�Z�4x�MΩ	�Z��� �i	���[R�en��s�EI�`_j11�l���\�j�p�_���'��H
yu�~-ڼJ�Wy��N,�\#ɦrYH��<$c� �I����P���у� Z.
՗:
��PIG��B9(�ܻ�60�O��Bƃ1n��w�1��#���X��K�4o����_�	F��Gă?�`<�c ��2r�#%Բg�m.��m�(�m�!��2ە��0�ؽ�}.�a<�O�:1�>sz8~��p����)�ri��z���S����X�)����zt�������)��xIc>� �$��?x(�����nr]�Ȩ�r��3��9���IhM�+t퀾�bت}���Z�kz��H�(e�?.��PMÖCu�����a+,��}Ey]v�+�[뒍��fv��}����qP��vYk�<�A�mv�稱F��n��⑉��N��x^�u�uO~\c��ӏ E{�Wy�㖶�ףa0��Eԁ����Ö_�Ba�c��΍��c)��F�Wm��:�w� �m<"�ѕ�k���~F9�-�΢�+ྗ@?K�V�y��#b�������D����LV&����ot�>����:�@��i�[����a⫁����uy�Jc��Q�������#��>[m��`��Fx���w�@��	1�����5���	�c�9q���T��E��ɫ�Fy�u��A����<]�T�d"[����5p� <��m��~[0�a	u2�������s��զ.�+�G�J_F�ňE��8JLzt�,Ψx�M�NAO�k:~nGvb��;���i4�NF/���b~��H��y@�-��)÷�yt��t�=��G�W;�ذkx��@-tG�o'O'N�N��:}�����2���:�����;|�w���n��4�x����Q���?�a,�I1��Gtx�֢����C����6-�p]�X��XXGet�8�����c��Ŏ�k���{���Y���3�����a�����q�Ìʓ��>���r�x��@}�aU��ac��?1�x�B����{�8��Z��{��l�?��t���¥��ً燓gϸ�h�YJYKq���'!���^��/�<F
;�Ȇq�qm�el ���D�0�_��Dī5M���AV]H�U96d0�d��ǅ�<֏�B��s����d����"0���~�p�~����5e��WF����#é2ʎ����~���5.B�՘�����Zn�Ǉ"�rk�8՝���U�V_���Ǌ���<���k��~裺�c���J����~v2�c�{7��a�T�9�>"�\���]OU��۸��Χ�q�8dT���T�v��|��������T{pa����AcD��������N�<�~ŝ�����F�D��+����e���ר#.�`��ϬS܉!w�����؉��ͨIbյ��!���2lŻ����M@�����ɇ�&�vcmw���`�.�x�z[[��]�X�nz�ϥ���ؗ��e!��f���������W�V����,���լ�u��D ؄��nT0�	�c�d1�2��i v|F͵�׀n��63��[�Vר�!������i�D5�b��:�;�k�ENYIs�/����l��
ꢖ:�%�4��݇����bK4�\l���;C?2lY,�IeQ=Χ5OhQ=�Eط�,��	-4,�ǎN�>����p�����ŋÅ����.�.\Ξ�0�9w^F���g�Se�j��@��Ͻ�v@�#�9�����ʎ�s{ʠ�:x�U

��>�"嗡��P+0�����D��A��'d��8�zm�g7�[�,�<��xd�_��~��*��OႲ]nȮr��鏊�����C�t,}����#=�b��n�F|y�#}(�GȈ�G76T�����ݯ��=(c��1�{���a��[�6n�C��|�����x��G;P��QwDE\��a�Q~�h.Xd�>�!U�_���s�mv%ڝ�J_T>2;��9*�c�����>��ʫ�"����Hs�B�Q/Չz�O9�w��%$seܶ���ؠ��CŹ������.�⢀�g.�~B�d����C�����e�R�Å�p�e����j�c�	�(V<Lۊ�^�!�)�?�)	�z�leh���. ?�(�wl��^���{��O�n������ҽ�x8x��plC}NF7�'xYr0��1��h�9�<�hΠ��O��:��+R6m Y�g��/���Å�л����Q������;1�v��Wƙn�@yUf���
=����+��v^��G���������X����eqt�>
�M%��jzd:?n�Q 3
��e	��d��{�ѿ������]/�f�0�Lu��$�H�V	�W�[&�Ӣ�)�^!�r�1��p�0j����E;��$������L|_^�������
���@V�V��h���,��v#�����r�g]���@����[q��y0���6�Q��%:�O���Қ��� �Ή�S�K�P��oL�ۢ�s{�8�ӋtA�f����-\�ϝΝ��*���]�	��2���w���ʥså��d̞���'O�O�6���(_��u���o�x���Kr��M>�yox��X�2G02���A��1Ϥ�����ˏ˟RhjF�ɽ2f1j��!��Ȍ������ath8uB2��٧�˷���L���2�x�������B>�ʷ���S�>�3���[I�Ez��B��+��~I���}����Xty��g`�z�y�;l#@�m]k�V{�+y��q�\��_u�v7rcW�WFn�x�%+׋/���RF���:ݸu{�w����gU��}Kj�K��b���ky+���pdjnr���r_�&T�bC.�%�ǳ���bj��¨�HܻG�&C���cÕ�燋���Ξ��w���:vA(.�x#2�G�_��V7U�۷�s�~��q������m�l�+[^�e�j��xӌ���-��(�q+�����v _��ot=Ξ=9�9uB�P�MF,_�������0p��.e�JJ��"߹wO��'�=] <W[���g�,�[�&P��&�j����I��ۂ���x�����/�����������~R��tAx��W�!��_����:5�>�L�q��pWua��@���nþ��d\�y@�+>��;5>g4����-6�O�k��ǰ������n��ЙJ 3"����'�adQ�<>�'9-B+k��ֱZ)���u� �mVD�)>�V�JQ��ez������s�V��4���]���9'ڢ�>e9����݌�2%���6Y��ϲ��}�2�B(�����46I���)g���G���jR���{�ǵ^��������oj Q �f�r0Na�0.׃��S3�N��r���f���~��Y���H珼e���"�e���O��|C��_�\��v�J�Ejz���hm�G�������SkԈi��B?�J�d��$�]���pU熊���攴N�$��2|���tiZB@����*d1����%@�����g����i���d8%&~!�~.#��O�?<�?jx�K���eH���A��������P�/� >sr8qℌB�CZ��sS�t�5XZ�x�_��E�3ܿ�Ȇ�W׮���S9���,֏��)�V���<��IJ�ۯ���;�V��n�i�s��9��~��Ŏ����$�~�^�Ui�[v�|�XF��w�4��9s���OӘݔ��D�S珆��"C��ӧO�=�E�Wj=�KF�c��㜨lBWL:n��ω�84�=�1�>�a]����L�<j�-�'x�Y���!v��֭w��9Ҹ��[�
�}�v�+�oܺ3\���p��]��E�[e�����MD/���������{�Q/�Q�%�J��T=&Dv�cW���ꂃ�?��ڃ?w�=��s���tp���������޹�c#̥�I�s����w�W�m�p�s��pK�����)�7�<��\�66T�q����/���U�~���3*�9�F:;�<��'e�ׅ�8��j��s�w�#Ǐ�M�˰�N�l����w�.��In��O���it�T"��k�ܺ;\W{�U{11�}Gd�xS���!�o��z��0�� �`uw#�?���;��E�<v�qlC���d��g?\pi���Nh��E�q.F�?s�$�c�{�s��E#.c�����ƭ[õ���h�KO\r"��?��.�U^}&���4���{,��u��xV�@�N^�X�u1�믙���?��Th�@�P��FԼ�� ��)�85&�CV�9��,K�`)\�:Ҋ_I'b]���������\2��n�pk��.�����O��zH]�8L O�镌[\ ������"�~/��b��T��5SF��`T��xU.�����"��i�'��l���+�d?�4֊4n����>da���:��`H����P�$ v�$T�
(Vy�!�<v ��hc�x�$ъ��_o��?x��_�'�nT�� �Eu�o
��R�I�Hc��p�������~����N���H0h�P0�),���h(��C�(�VQg�@5���GZPQ`p<1�G@�b~04��敃N'�_�^�K���E�"��Ө��A����w3^��ڏ8���z��$��Ϟ<�´w�x����;W�����wߒ�{~8����]�����Vn'�Sx��Q/l�ǂ�d�?��l0e�L�细�2�h��y��p�����}1<z�І�ŋ�>���k8w��w�0n�<yn^�
1�׋*Į;�'$�+���{[|��~��p�������{�����q��q@2�ۄA�{I1d�����?��ʈ���[������S�������^�E��2�/�H;.����Xzx��ϼ��F3cӓ㙹�v���-�$�0�<ut�D[�}I|/�/�d4k��
��r�綱�}2t���n�*v�yv�
^_���l�_�qs���W�_~)C��z��`��6�r���ᜟ�>r�����㮗�)�P��T}�>w���k���ᇀ�lJ��2d�{�w.Kw�U���ϪҮ�M&rW9&�w.L6d0a��q���mo>ٌ�.k�wOR_}}s������o�l��Ɖ�*�Փ�vAF�I�9(��+)/:��ԍr��q˟�Q1�����������~��.�2��70�y��]\����C6ԏ�,-4�;�s�o���ت�����Y��q��}���>S{��͙�g����E��ݑ���a���Q���CH;���Vq�_��Q���!<;~����9����ʥK�X;%�����=�����1~T.��y$�9 V�_ r�@�g��#>ǥ�JgŢ�U����w\����qAs ����;�/4g�˪�\$�TU�1
�x����磝�ͤ8�2jð=Ӕ���ͮt�!D�:a�[H9Y��L�ۇC���A|�p���U�˂w\ֱ���t"�eR��/7����C�n�����^���S��1��ԧ�6��j�wY��v��϶��p�vs��/r�O�5����Mo�a�CYZ>0� {���/Ӏ�����L�G�.���O~U���;D̍a����sn���D��tU�
�Z�Q�Ra���� ��Ju�Q)��/�	�1����[œǊ�r( +<4����h�i�a� ������"t��E�Z2n�R"q8jj��>�5��7��A �c��q�T��~x�IXg"�ψ��/�	��Z�l�K��2p�#�����)��_�Ƃ�RA�ծ�Ff�2�O���y��9-���wY�ۙ�̩c�A�e��z�ƍas��a�yFu�sDB����~�X�w��w57eH<��x~��v���nٸ�j���O͛�߫W.?�����d����-�;wy��G��cD�\a����� ?urcx��+��޻*��p��i-�G��ݼ��;��Od 풡�N��}�mP�Xģ܉���2��w��Q��U�c�2Rd�>{�r�|����G��}������+60�x����{ޥƨgj䝢���n#���2}���p��������ի�o�=.�`>�?!�s�)Y�˰a��%�^�q�v�>��Ç�Y/⸏�@�QxG��.����7d0]W�({�������/.\8����C�ȸ��m�ؔ�1Wy�U;�(���^�ː��	y7��S�d���xL�<?��謁�åK�l�p�X}��[����c�zM%\�?}���0ڽc���<m�c$������-?�@<w�Ȉ��8���{�ِ�쐾t{�S���W3xl�ʑao�xb���ɣ��:/�qQ�Q��(�j^ѵ��2=�c���.�7��Ý�g�CoQ��k�x��ꮱ�c"�'񎭌�/��j����}�u��I�{Y}���������ޝ~���Hc���E]XS0n�*ÖG?xl�.^:k�i�˗.������u���˗�@�����e��9u�;��k�� ~&Y���}�O~L��A��]��E����m�޸yCt�U���Ug/����K�x�L��m1h3i������Ys�F*<��Ѩe�KÖj3�G��XB�����ڐ������&y8O��X�,%G�n�XU�J:�2Mb�?��.=D�)�!1���M٣�e���q Y�S��g��@ұg�N��'L���2Q��w�&RJ��ܜ}H)�q� �g^�㼁$)0+x��#�J����)= /cʈ}'Z�0�ܑ�q��Ӹ� Uc��Xz��oP��_�R<�� h�*b"�����������(��rU->6H��D/Wt�J��P6~�4SаЧl���P♾����x��F�xL�J���.>jY�� A�
�)�(<#���W$�2&�Z�ׁ����g����bT�5��`l������p0��8b��D��g�Qb����3�[WN�N��-���p��=����_}�����ݏQ�)��p��3��Bxs�q��p��-�ݱQ����}������������o~�w`�:%cN���=���,`_^�=ܼ��2^����#���3p������}����C�m����'��F��uu�M��Q~L���a�����/�_j��B����2�o��چ;�{��L'���{�e<��w�����/��-觇��Ò}���>��+��%C����g���i������g����Kg�w߾4����H/gNm�߫�������1�t�y[%����=y�Ńt�����׿�E�����dTܖqw����sG7o�	T[��®�����|O;��>&��E}>��6�'}��-���b��u�ƻR5W��N4��9<zxW�K�ٹ�����>�������Ӫ�~��h�Uvoy,<�-&t�x�������6�	�[��ta$�:~�����	�<6s����O��|���q��Q���Ƨ�����T�TiՊ��^\pџv٘}KF�������sgOJ��2Z��%��{���<������K|��|��>2z��6c����-�,�~Ȏ�W_}-����Ͽ�q����_L���.dܞ=sN|�"#��ʎ?���#aܪ}�Fğu��?�=V��O�E�o��.l6�S�}�q�d�Z��ؐA�D����/\$�t�;�<����ysB�u�B����_|9��Ï�k���x�N�{�{ox����=/�v�ރ�^H'�'��ߨu�{t�0ns�}��,~��V�ؠz��/�Ѧ���@[�`�鱠�{^3��^���cO�;`�d]�j,rD�˴sؖ�G�.�>�q��cʖ���e�3��O�r�W6n�6��Get��E�:����H��H�$^�^���|T�|���>2&=���L��Ђ���F�����$�̭.�Oj��0&*�X�5d4������j��;b�Y�o�F�|�d�`�B+~��/��?�3:��6:����3u���Hx&�<�aP���y�(W>�`�v�:�c�C������&��u���j;�T_u1��d�]P��<p`��}�xOg`��Yt��iEcq������}���W�����_�R�_�~򛏆�?�t�~����Ǐ�:χZkU��Rt@�=��1i<�ȳ��G��G�}�������X��W���N�2��w�A��UC2HUP��?�T��5��<��dHݖ!��_�~�����_~���ï��2�1�ib�?�O��?{z8w洟��yX���2.��TƮd?v��(��@��? ��&���i_d�h�����v���'��N�:��y���(L�1���q�P�G�DƎ3�2������eP\��.N�ې�#C�]u��qH�҅
��������9=\�tJF~�P��x�Y%�d�]Ұ/�9a�Г:���4ء�c"2Zy^�?']8wR�i�yr8���ĳ�d�S}D����+�n�H�裏�_��WÇ�f���O�������O>I�S���1ޱ*�|��?���	��dT]P[^�xn�z��p�B��Ʊc�%5�Z����hK�ݒ1C�.��n����u�u�sq�#2���w�����ǟ�}�y�.�>������/�u�����=z(c��]��/bL�9sB���}�>���ct2W��D���k o(��� �Q��/�S;\8/���ѣ�.��[����}]�r��.�낊; �7$+L�n��Jc�tvi��x(�y�[M��Ϟ=��(빤��{t���1��h��7��݈~f-R'�HbT.�@�1�<*>��?�b+��0��?�� �U�@x��v&3��]�~��U�[f�_��u���r��$��@Ӏ������<Qi�X��BO�����&_��q���˟�����>x��,1���w����3�>�k��	vP����`x�J�;��J��y��w�X�@��УQ[�mM����ǫ��^I���:�G�Э���6�x��./�,J<�x��>�=���1���ڟ��� 8@ǿO�����_
%��CV��n|5<�G�Q�`�oknk�8��U��d����
6�Xl��c<ԟ?@ab��
3�#��V�/.���k��%:w��p����s~�g
w�����»��7 <�ޞz��8rX�q�A�ҥ�Õ��s�3�i�dL�ox�րAkܣz`T�Pt�v��!�FҕX���^�T6F�8�3�BޯJ�<{��R�;=\�xYFȅ�ԉS�@8,ֻm�޻{�/,׏�<��>~��ɘٿ8uZF��sa;�E�u��{�CEb�S'�%���O���(j�~�p�d�,�����3]0�7�4�M_u������QR��o��W�	��\�����f��=��W�����4t?�TƢ.Nx���a��W����tNmN}�������{�0���@�iP�g�}�O?�]W��P����s��:����S�u�0��#}lc���������O�	we|���/��6\~u�+�_���wl���;\`�����
��w<�q��(۟��P���S�.zx��5bN�[�J�ng��31Ĺsp?����ݺА�G�KG���Pe��ϩ?�l_^�6|"����?�P�����g��g�ǺP����7�f�B�ܽ�Rt!pXm����ua!���eK.>A��D�q�}.>dA|�q�%���2nuRMcNs�̾�<C�T�Ϲ����5���%Xﴄ��c]U2^���׵;,����B��"r�?62V�,&=�U�Yx5n��`(�G��E�� �*h�0�4�`�'yu΁�����%�"����}|蒉/&���pu�����*j	Gg�wt�g.!��V��d�a����o�C��U��a�c@��(]��c"jx� ��yĸ��"���+�/�=�0*��$��0�Ta�͍����?�y�h�֜vދZ����8����S䵌��E�<��F-�9�g n+ǛJ�5�D���>І����I��6/K�˗.�e�=sF�����2�Ni�=�8ˈ!,�<���?�`��<�1=�"��t%����&N�oDr�j�6IS�0�=�a�SweF����1^bQ��;y��p^��9sNq�e���:罩���~��É�'U?�qN��(��'��J\�����S��>�];�"˗�����'&m�<QO��0R�"W2>hq���
�4l1L���-�<���xV�Wd�(���(�-�y���S!�Cmz���᭷��\��v�Ok�J,�f�R�� �m���}6:����D��ꊛ�֣_��-�t ���:ほJ�a�[ Μ:�>wix��[�{���Y/�5.�(N�Ō׹�� �rV����.�iՋ�	\lr��+x�m���@�}o�Pڀ���D�p�0
���'K���D��z<~�OG%/��g]�U�x��w`g�]�k2r?���Q̏�(�]��n�}���/4xU V|��w�W�^�|��0X-��x_o�2.@w-��8,�Z�́ه��Hr�m�9:p�߮�	̂o
b<�����-�m�4\����9D}��R�+@�'ƭ�S�폱7�	�4c��A���1^{�������g��y[)ɋ��bUX)='m���(XLpL�L�%��p�H⁙H�|��Ir�[ �F��O6��bb~5x)dɉ׫��5#�E�%�l�!E'�HwV���O�D`F�a]<PY��YH�lL�
#���"��C�B��M6[
�:B�a��.W�k;[�4�{���w�:��'0ڱ�,#<YD�c��w�>���o=r��������Ν�����������?z��Z�����uL|�aC�)�GRg��.\�Z �]�8��U�`�w�~-x'�SZ�����f/�n��=~�ɍ�˯���<�"�\}Z���O?��G���rz�����By�o`׍gu�����4d�ɸ�4����������p��i^Ʈ��q18->��Z��+W�垻xi8���G�dL��w@:{1�Q�2\؍��ӧ�������~{��Sn�����1ʹe,ͻ�򶃽�#��ܼ'�t�.�x8'#���Z����p�����׷��k�~�{�����^�Oī�x} :"��ĉ�n^O�1u���z�dh�q�.iW^�ϔ��+0`�������|�y����_?��/�[�����#�Z=G���{��0�����y���2������{c��P?+��ǟ�uW<��?���������{����7�;��/�O�>��ˎ�K?{�wd�^U�^�?s����3Ȏ!.;Ӽ����~��S��C߭��My���q��e��$�+g�שS�t��+�.��7U�J������`����ҏ~����t!r���0������-F o��v��[8.^Q�Ϋ�ox��
�����b���޻�\��~�돇��Ox[�}�ƴ���,�G�hp���O���H�[N��jG���q��tN�>�:^u=.Iw<��L�����(b�~^'|��r�u��E�O]��m��8>�:�R����{���p��?�\S�wŗ?[�E󖇎$cn��H��n6s?����>~"�YtEO��wЇ`1?
�,�S�����,���y>��N��+�9��֮C��X�E΀�u�vkD�C���꧎���qF_�1_���ZT�w�̭�́,�l����8Z'�^��X��.i�YZ�*�1eqy�S艣����c]���#k����<W ��CpB�bj�N�Gy*�C��,?�3ES�?���:������Ԙ���%�h�$W��7�%��F/�V$.�ڭjǅ�5`�)aj�3^I�
A���R�D�Q�'���T�|�^�``�N����:.!n<��N�AV}̓胸`hb�<�"�G�8��]�Q�k�d4��(�<\}��w?�}����w�'�����dj��{��U���_N�;?��ЕyEF��o'O�񫂸X�x#P_��ڋ4�ڳ㍅z���(��N�o�����O�����ϯʰ�x鲍�2�m�Ax�_P���;�;�{x��0\}����.�4l���G��� ���nh����-����IK3z�q$�Ƒ��g��a��ˀ�s@q�U?	��.���N��j��;���C1�x_�Qɂ/\�}��S}ޑ��wU���K2�/��.^�<��tAgeT���L�
;g��+������-*�N�&TvU���Qm����c�����0�h��2�'8Ȣp<*��$^X&�d�������=�/c�?����~8��6�����~���ڕ���"w�\Dq�tZu=#��J�S��C���c�͡�J�!��S��;�yg�.fl�f;��]/��H^���|9�O�����y.�p1����\h���a|\6Dwd�\>c-Z����ʗ�Ϋ��4��^����Յ]m��ѫ-%�=.,o�۽�5n��EV"��c|$A�/�R����/� ���c������`�ʅ�tF�I]��Gv�VL�[F����Ǥo>�}R��\o��p��+Å��6���<�1A���0vy\���s�U���s<^�c��s�`�(��#���q�l�;҄����*�w8��3��Ӓ���a����<9���ȭa!�N��2��D��N�>��w�?ש 2D}�s�#��^�q2f[%6ҺO��S���?�L6!�_&�����@����<qW�9�"t$�����i���*�c���U�������<8�C �x� �JN�E(�˨���0�h��q+�E��_W9�ؗ�{���s��ʹ�DU�*(��[�NI� J��fB�V�ȯ��Nlqԙ�wQ�`����r�s���.�![�\e��E\wd�(����$�b:�,��o)��7�HZ�1�'��0%TP�~���S��\�mқI��ˑ��Gz��3d��A5����xY��c��>���O��������G��φ���������p����po8�-�Wd�^��}J�����c2��Ȑ<��4Xn��8������x���b�jQfg�Ŵ�_�����"�?|��$OȘ����2�޳�Wr?G��K���>+B����s����pD��c'�}��_�+��Vl?�������]�X�o��%��Ƞ�w���Jn\ɊQ����a�ad���E���U~y�.����n�ŗ�QƆ?�*c�Lh��Q��(#�n}�{2�d�^��wAF�H�ϟ6d(���Y^^�g��ʌG"bΈq�81lA��gyc,�H�'_7E���S���e{���e)�3�KS��y����G|]n�/*Hg�O�޷��ޏ���<������G��zKm|Y��.NԷNȘگ|b+����y3�-w�7��ȝ�u }�ۉa�W���y���R.��
�F`��Vy١=y���ԅ��2$%�E� ���￧��k,\�+������� <*�������7V�G<�zR%<��|�L"m˕n��0��:���2�{0�]Ƌd��ާ��1H��T��y��G��7�ʃ޿����{΅�������"��;����|�#�U]$B��N�9%cWc��<t�\��U_��>���L[0w�7��/U��cL���M�T�5����G���M?c�N�>�6
�L�9-�R�i��{Ǩ�<Y�r��ʅB�}�M�nG�/(��X�=MA�M5��H�2�V�����K�-qkX-�GPE�s��GwJ�2:a�O����:^tЃ�θd�h	��`�c=�Bͯx�g�͈/��k�JH��nw��f��@��I_�C��Tt�?諅%C�N��yv)�*F��p}�����s\�V���w��߹��s�6$���Wy:ԩ�M�ΏRR9u8y���8%GA�	|h@��Q��xų��8{x���ʗ�ׂ�u
n=����QNHK�ht��ݹC:K֍�_+Y�B/�ϒ3K�Zť��W!ˍ)�Ǵ�'g9M���d��Yu2��Pi��6Isk�6�NZj3#����Su	7��5İc�f�g���2/]����x���ŷ�3�.'O_6N�P�A{��qsG��^��,b��ܭ�Hn����n�G�~Q�Q_`� ;L�.�o1k��L�BW�_�f=�!��ر(#:���}2ِ��{1h��(������;\R����O4ޭ�L�1e�i?�i1Vv-o\��a��k-�����2�0~cg�6v����l�*�6��x�R<gJ}d Ȉ9*���fv �<*C�t}H:8 �b;�*��t���eR�/��ݲR����%2iZ��EK?�1�p���J��ba)BՕz���<FFy�jkޛz��q]h����f^�t�;�ܶ?������3�\ȳ��I��f�� �V��D�:Q��٘���Q�?´��}O���N��l�A�\0짟����ٰߨ�^wG�N�t�!cQc��A���~���!(�񜯿D���~oU�:ݧuUbz.���g��0l�H�����ȥ��m�᙮��<�tA�8>��.,��;|f�w{�ˈ�����)�;ϧ�^�ݚs�y��ف�j����}o"}��[r��*S}�k�ɘ��鷼~����4�Ŝ/H� _r�^h���6�99�@��M�� 49$oK4)���e�)V)�o�;��=�aS�I�q{s����1t��F��Mf`��W��J0��$h^�\�L�������p	��%�u,���F�:1҇���uѸ rj-3.WIeQL
�������� V�թ��>l���00�g+��w�ɺ���$A9� �:��ξ��MC5��-�R%��A7r"�S�eQ%�9V�[�1�/?������G�W�jjQ:(�ވV���#2��߮<�t�aW��Ö�:��N��l��<'H���Gx�5>
�3p���k"�$+c����2a<)���0f�k�|*尯�R�T<�J���"��_n�b8��X{wՆd������,[-�Ih?c�� #:�\�k_F"� �2��A��Z�7��/�}��~���B�%�Ig����[��je�u2�l�J��̏?��-�Y�ّ��]�	�E��Ż�2Оj�x�����M!��D2=1�z�20^���R�w���0ڕx�K:0"�����J����j?oRr�NYѫ:p���|�P a�Ω,d���n���_�/p�Sh�3�>r\�:�!<�>���Њ�����cq��
�_]�tЗo�C..N�/������ݥL> ���i�	�A�.r� ����7e������ɳgd�6tarhc�;�<~��.����G�yU�����e�BI<�ʸ���_i:�.��i�+Q�n��ry���~�c���2ry���p�
;纸�{������82�gHZ��/��l0_!|j���\�U�`�a�\��y��y|��oI��7��0���<�XO>T�"q�W�| n�u\r�s@�ܧ|-�����J�����A_��dS��έ�%qM�C3����PGS^�[�fU�;���|pFw-��'��+�����XqS&=�i�j�z�x��2��T�Z#,A�oAX,t�[�Gdp�X�c���g�1ț�;f� �B��i{t޵ MLb�G�U 2�^A�KL�.�O�NA>�[�<�)Hz�q�:��w ��$Gō�1bL��)�w�2�ҙ�M��K�A<�H��H�~�m�l�E�UvN��k�������7�k_���{$�������އ�2"dY=y�K�-M�Q��q��p�ƽ���w�/���
�n߻'�C�.��c4��x�OB�!K؟�U 0+#a��^��.d1~��x�u����������GO$���(���ӽ���p���p��#����񾿎��T����[Snx�,�2��W��h�u��σv@���^�����Ű{$������]�xW� �����d> U���y(�#��\�{_4|����~��}>�,��:�1�/����K2�qԸ�}3��V}�!=L���g.��W�,��84�S���������P��?>�a;�}�A{޹�p�u���H]i7�ّ��YzB��aTX?t;��lw�(�����ݠ;?v&�һ���.�������0_L�"��U%8t��G>�%]JV�?�����W]���b�;��o����[\�[W��cշ@��(���냛�8�~�G�gW�8!��]�eԞ8������χm\�F��j�1+��y�L�(�zF'���Ȋ\�a�1[�-��`0?�	��g��ׂ���cM
�p�WkM�߸�B�>�DY���F98����g��ƨ���u����N6'�.���S�YI8�i�ׅ?�W��-�\�C�AT��	Sy)���^؛!�z`�Y�%���p���LX��0s�}��C]�No�^;�u6q��r�0��G�'`v����	o��fr�Z+:����nףH�9P?�΅��l�� 0qx���qj��b�]�,� :��P�����'o��������}Z��G�Ч�|>�짿~��d��,���P��}����u>
�Q����_�������~��φ��������G��������p���χ[w���-���l��K���^�~u(��<��e;�Z|�0���~��g�ǟ�ڢ���7�7�� ��}K�m@�#���y[��M!����D�xu׆�i�vb'Ozd�7@�Oo�G�ѧ�'h�IP�T��z�1�M�E_�5�r?�N��9^�F��]������X��7��Ah��+�ƭ������r�^7��}����g__}��pWm�]$m�'���N0N�������SȄ���M�/r �籄��[\P�}yw�B��s��t�t���:ݢ��ݮ�n_��}�/z]w$L���}���$�؈��
�r�A�W-������Wڈ��,^���gٕ�c�O�P����=�"���� ����V/�_�eP�Ӆ�]���.�+�N��"k���w:�؉����p�1�W�-�ɂw`�9`�i�k}ܹ��	_P�_sA��<2r�wn��@�v�;$����*�d~�z>�K{�0��P�2�yn�x�-b���n��z 1��擼<w�Nm���$�L��A;��L`��Әv;���<*C������0g�����C�W��7�~��ۣNJ����!�"-~�o	}YQk��g�e�z��#f[��S~3���2��U���e����?���@W�H�z	_�4���K��:9�W�H�F�*�.:4�a��PC{�Y�5�p��A���;^R�_�Ţ$�l)�=(Z	�Oy=���٢3Z��H����`#\��$`�8A�˲�Ot�8 S�
��Mx����\Ѻ�dYQtԯ�f(���3�[�C�=.A�'*܉�w�\��p� ����j��'�g�lΟ6��&��X,��Ⳬ����W�����4�c��>���~������~�%��g����|�H(AsC�7�H�k���,o$دzP��ï����O���a�����hA|>�e-^��gCO�>>�'Cvk7e�ܽ_�{�����C��O�x�fG��Kvs��_U��|��֝�,-��-�y[����B���$c�Wh�G�c�������2J_��	��ç�^�~��ϲ���f�\�gz����������~�,�B��`'���P�~�A�n���ãǛ202����T}������Z����2�ϲޕAE�����=��/G��{/_��/u�_67e\�z(���O�k��n�&����>~.��|x��?;r����wn�e�����U^v������k2d��
�nC�?e��*;�|7e��3��X�b��wy�ݳ	�m����s1�X�"�#�8w��f@�>��9|q�⯽C�n�SE!t\�}�/���d8��pb�_��_�z���q����<V����|Ջz]��߾)����S�I�;��zܑܷ憎�YkՃ�����xo�ָ9�C;��*�P����>�����w��]�׀1Y���s�V���cU�m�O=N?��R_f����p�Ye�Z��~�����̥0��*�ݽ���X ;���?�I/���pϟ%~�?G���Ə�q�;Ç~�y�g"�l��0f��U;��N4s]�w������p�W��T��sc����f�,�a�	<~�
��4?y]�� ��#�9�8��)�
T���������Z��y8�䱰��=C�}8h̃���e�&�#�/(L^|3'~%�E�w��@"�i�(��o�����}��������}��������E<B�L�ǬDc�:�Q��⤢���$3��U`^��N�<6�y���G�����LK��9J�u�-X�o�[ezp�BIs��JP~n��'���4���|P��6���&
�W��KcΫT��]?�������,lZD"@Z��ô#6�5 r��P�� ��|� I�!e������Y��Sn����e�?���B�>���JFά3@�� r�QSZ��ЇI(O���n�ᙌ��Z��S�ϟ��U�u,�}+���Z��h{ ��wB?�q���?>�DF�g������/�8]���g9���ڟ�Ԃ�|��ܲ����}n'NĿ�O�8�ҳ�ݔq��G|��g��1n$?F�������#�mܾ��U����2!a�b0 '���[2&d��P���/�ϝ~���_�Vx�+9�",��W��R�/��/>�[�����!0�0ny� ;nw�=��a�V����'�
g�`Ǉ�v�����sO00�W�._<;\�tʟ!f(ߗ�;L��q����d��?�`����Y�M_��/u ̮��B퀑�q�'R���gn��d�_���{G��Ņ���U�
��7o=R�~5���ʸ����m��	s,+�g����[���d��q��}�P��~�-}C�x��K��Mߺip��� u���	X.P�P�Pĸ��>}�T"�E�#�t���˕q{�������2ne8sA�ZqR�����H�'�_O4˸�y귗.��y���s�Bv��!�χn���՗�ǟ~,��_���}�����/�O?WL�_�$�'�m��S�u����S����u|���˽�Eƭ��H$4o�Oe<����}h�����-���:~د`c�~��j�/��zW:����������ܽ�+��/�>ׅw��R�Omr���5�i�3>������;��|!�ڃq����yb^��S��{2�^��vM5�bݢ��Ě���� Iv�'�%;A�T�����shB3lk����t<H(�K��<�Z�������;�:g=g@ѵ���q��0�"�#��g�
���B�e�/�{�����fj���?l�>�a���)M��"��8���ĸe2p�H��I.o�(��!�(�x0��U�1t:* �ę�d�θM���C�|tT#�=8��E�r�Pn�Ҁ=_�&lzZ J�3�I���(���K���l�LG�D5���W��c;����X*˹Xn;@ʔ4�7}��N�w,�
��*;�on�Y�%Xv����-H~��G9�2�r�P�!�>J�F3b�m5-���{ʿ����v�XH�<ת�xqݽ��R�ӵ|B��Cþ���������p������{�C[�����'2b�J�ӧ�§�Ƨ�g���L<�D�PE�k�{��LC-���ؕk:+�����q�=� ��?h�k�xL�.��d7C��/(ݔ���z[�{wdaq�XH���F���1�&4�W�Lm�(s2"�(Tח���/�#����<�� c��U2��t�����<�1j1>0v0�m�X���n�H��e8a���t��w�����W��	_��2��g����$��w�:	��lȨW*G�F�g���H���FS㢁�r_}��J_ʀ�X��'���XB]D}-����w.�h�{�E�S�1�rQ6�'2Fm'� ��0��B��F��ދ0�����x_�~]�g�D0mB;�F����	�_����|�ߤ1���G����r��EwPxK�EQy#R>u� c^�~%��`�c���f��j=���w<0H���?���7������_����/���r9���(�o1���	���
'��/�*N��*����P,����s��1L"G;x�h�R�6f��Z��-#3Z"��|G��~����*��n���D T��t�+tVy�p�^��Z �n����vVu��a)����p.��B���pN:2݆8:�C�j}�/`]aE����R��)Cb�e�4���0aCY�N ���4���:��О��D�+�UE$Pcb��W�5m8%���y�)ƴcC�9�T{�I�,7wi]>i�s�Q�G�R|n�Ey5�G���KPrP?�u@Y��,��).C�o�/�D��,��Z�e^KP��b��c����1�6^D��j`P�N�ӪE�����'�5YLA�g%ge�f��7¸}l���vǷ��7,�Ӎ����G-A85\�rqx�ݫ�{�{{����>���?xo���w�
+���m|�+��o]�\9�m]�t�_��v��g��ù�|A��p��р���0�"�HV¼p��:>�������wX�`a\�N��ďg��9�Ϳ�ֻ�[o�3\�t�/�?y��p����TÓ�ϧFO�99�9wz8#��+d|��ԩ�_k⽩|��Б��>]A�F|4������q�燹��A%#����g2J��Wƽ��m�c�{�7��#����ĝ&>"q��}<��;Si+P��o����aSț-0\yN��!���G~��C]�p��T��~��׹�<�k:s��(�_��2⏑�����6��t57X�%�r��P����B������.?[ʟ�h@œ�v��Ttz���/p�>{J�C�t1��P\$=�Tuf|n}��ş���'c��S�>������Z1m�7�p�=������B�b�T}+��m�\+l�z���|j�'/����x4����[����7�m	�x�Ǧw�ٵƿ���}�C��S�ю���m�����] :�?j�ϣ�K��6���[�g�'h/��ׯS}�x�����2�?~!�o����_���
��F����W��~������k��?���nǳ�����~���^<���X��w���-�.�'���[�+S���[QP�W�窛Q�:r��Q稷�R��˟n��c���9t$L���w伸v~!Sx��
*�N`\w� ��5�.��"���F�*S���:���נX6�xP���#����(�N�S^ң=�V�1�m��]���~������Q?֕��Dy�?���y�L��?����s��)�r��q�W�J(�T�d�D'*
Ax�ڽ*TL��ɝ��&0��������x�C|���L/EQ�� �\��	�hXL���q"�D��k�8���	ހר�
v��n�BEp�:0�B��"W�Em���zL袂�e�b���p�t���
�C�٤�:�V�S�Vv��-�iՆ�QK.�F��oB��ӹΗHz&��Gm0x$��w��A��?�0���1=�Q~����q�K�������ge�9�����������W�Nn������aH�i���X4=_ʒ�H����"����5����v�%�������e?|���>���9�1ʗ��#I������^>W겍�B���U��J�w��N�sFu��=-��V����o?��~g����3�mڳ�1m�\����<��)�ȡ��[W/��. �GT7��lQ�3�:|x��W��X|e��ȼ�/�m�/v?���ЅD|�u�.�@=Ν;#��W9�ũ3��Z|�l�A�t�~�K��O=�Y�CG6�X�m��fa��U�>�,
���geЩ�6e�>��r��p��������gnE�:�S�.�اx�ot����	޵}*��vL��q2���?�)^�4��_H���y�;O�����Ϳ�t!�t���g_���v�ό��_2�y5�e��$#��a���铒	�����<��7]�Ȩ|�u&��.Lx���\�N���v�v"�g��݆�s��pD!|Z��J?�������R�ڭ�y�~���_7o�U�ӘQ�洃/���%w���Ux��_�y����=��xp�����ԃ�>���G�}��$�>�1v�X��s����~^�&����.��b�]y�5����9b>��E �%���vG��?_���~��a�01p��r~����4`��{��g:���������� �؍����������o��%5�����Q�.nKH�	�N"�BDS:j�<²c*:�#�R&xb��c��j1��@�'���ּ���D ��C�<.l�����$AcFy>�W�q9�	{�qm۟�A��o ��Z�1�Jϼя��2 s֝����j�u�θ�7<���������䟶w��l��������򩐮����]92!�k*�ۃ���1�kkD��K�q��K���q{R~��X�w'J]A3@����w�T�*lq��mPW��^���om��%�|E��F�J�,4���t�̟���Fz��	ĝ�¥���i>!�I�=t��	�?��)�s�{%���<�gH9�j��e�2��Jg�Q�o)�y�|��#8��w�ȫ��I��St�40[ڃ�/tr�%���$c�`�`Y��{Q��i�?\s �J�JѠx��]��y��g�p����~����?~o�G���pY��l1ޟ�~��U^/�N��E��t�'��+1� �n�eW��$HT�U��/�����,��X�/?�>������ןj���C�~K Fe๣�wo��?��}t�������'Ï߿2�<�G�x/��6�`<;�XKNe�^�/�,�O���c=L�v�ݹ�#V<�r�}瑌���O���o��/��>�6�G^鴟/��`cҎv��P.��������k2��������'������% �(�;X�2�y�ԝ��^a�j����ACt�#� .N�b%�ԾbL����2D0@x����?�z�����������9���k�0�A[���j�P�"�̭�R��߽�Ű���p�����?�'�7��?�}����}��;
�#�#�$�nw<#K�ԅ~
d��Qj�N�ˬ�%�ЁT��������CÉ#��C����'?����o���ÿ��O����_�n����<�C�yU�����Ӈb����d8%��ݷ.j�3����`�r��o��Yu֚[���^~����!}�ƈ�Fvޒ�,���n�^;�Ѹ�.z���)�G��G�?�>����W����?!�������ʽg8(���'�?����3�!��勇��o������?��������8vXtj����h�%#���VYcG�Nɤ�$ݰs����O���<�Б��վ�+w/�k|�8~P�����[�}�B�1l?��d����h�W��;���J��U̇���J�y�B���;86pѤ�e�\n���L�p��}�3�;��5(O�g��$�":�d6��A\N�)=+/ʔaQv@љ�yP��c����y��Y`��"]��>���xjR�O]��[��Ǻ��?PR>L@��!���&�k��	�k�d���� ���/� Ɔ+�1���O���y_s=w�b��Wr���8�t8���<�˝?�8Fr�3�N ���>���xɜ'd���*��=yt_���l8s���w/������������L2�b�A�
��[8��RInD�tE�q�����1n�f��x�e�$' �@���qK'G���f��'�0-��"WSG㖎��u�	���J���B�ƭFb���Jﴽ��]�øe�ǸUٴ�-OzG��`�1���p�"=<d��ϟ~�w�ߗ������p��)-�2<\Y���:��c^z��Tk�;wQ%����V�kj�Q'�B[tS^1�q�����N�F���*v?�Xka����ߖ,φ�'?������ٟ?�����	�
����&�� 0qÃ�E8�=Q�F����냂U�������~����k��9iSu�|��$?��'Pd�~6<~po�w��pN��?�g?��O~0�ޏ�����M�(#M���fO�>�
����Q$'�x�#��}��͍�e�~5�������_����W��c'�]�6�ӸD��*M�ƭ�w�����棻�-�'�F��'?~����'8�}��.rb"�kb���� #�?XZ���C>�ڒX��m��|�z����}���������˸�b����l���>��1�R�C�Z*��.͓/x���c�קÙ�Z\޹<���;�ٟ} ����@ t��C�-eK;�B�#"B �E�?r�E�\(��h�@�9tp�.L��w�?~���������o�z���0n�k�?�{sY�PV"±ɸ�5l�uz�����z�}����#���\n޼�|��[�-��uÚV��My�B��c��n����J>�B���ޅ?x�u���g_>�ݿ�p����n��/0n��j��]Ɏ�B�/�A0e�+ވs"�s�	zBB\��p�9m'`z���_A�o�Ay*_�1��7�9B��������KFC��Х��yEkz����M��-���'���E�:�����k�Ը{#ƭ�^w4�w˸����'q�ʢ>Y�-�5�1Je��3n%�;����C4a7��+;����$$�-6��q��gߞ��ʸ��mF�Q���wgg*�IqLN�_���i�puJ����Υ�&FNF�(
c&Z���E٣��������D�W������kU��E�=�|�IPUĭ�	��TD�{%�qBOZ�4�5(w�N�]a_�|0|����/7o?�<x9�{�r���4����|�CT�߈��B�kNиN���s��q�$����p�ދ����õ����"x����ݚ�vO?�a�dD�X0���w��9�����cK>&��?���(%�4��l�T<g7"�����(Ѩ�F���(K����T��)�$#Z�=�E�W���n>�  @߿���g+�g��q΄ɝv���4ܾ�x�s���	;��Ke���n��D�<|H����N�/Z���$��R'*�Z�s����6��<�q��@>��O��h�t3CPy\+2�S�ż�)�!�~���}o�����X��0	���W Ȯ/�_x@u�P�4T��e�ʰe�@2t������o�}:ܼ�k��K�O�v<����z?�9؇�G������!�Ԣ%���QWD�Lc��Ȉ��=>�Aǳ��ÁG��W���A��7n; <$<8�8跙�<qh8��9�G�S{2Wb�r'Nr��A�Z��b��%�+�,�+�ƅ�1��h� O8}zc�p�ǎ�g�l�=�Gf._>9\�zJ������ꕣ�#�ի�_=���AsI����*��qϧEwf�t��pZ��v�Ir��?;��(e��Њ����ɲ��kj�Z�H8�|�E�h�Jk�|=����W��'p�	�����I�צ)���~C�Gz�>���E쎵 :��+���1��E�Q�^.���/���痼d�׾��^;1�H����[K��[�(��;�p��έ�5-?e��[!��P�~I=,,����3vmue?`�s��z��W�PF��sEPK{����n�s�$'DZ��k��= ��[v�r���z�"zP��b"y1j�1�n���_�)(�+D�o_aT����e���έR�S;��z���R.'P��vR"�@�PE7I�U��!M�M߭��\��]�; s���2�#N�
���å�� ���sq�p�����3=�F�.���k�	&�,n�E$97k�s�C���S�Nz!�UCC���O��>�1��_�j��ӯe`񧠸X!ܒT��cu��6�.]<9����޹z~8ubC�rW�B�yh+e�~􋶗+P�eZ�H��@P'x�:�(�p�|�k�tq�ٍ�c��ч�����^���?�Iv?� ^������c����|����.o�}NF���O^�U>?��r}�� a5#с���(�-�z���G/�k��_6��g���q����m�d2���4�t9	��&V���x�a���{í�ˈ�3��Go������,C�ڑy�qI�Z$󲺅m>"�"ZiAC_$ą��� ��Y^<�A
��(��o�n�"�Ïn��/>~�/�/��5�Vw|�l������{5nvOe@>��ydx��K����;�?����߂�0�A��p��eWG���|��>�T9���&�F��*��I�T}����n��χ��k��u] �';U�[3���VoA>\�I�Ë��e��������{�ߏ�E[����Q,[��US,@�+�Z
���}W�ҩk;���UD���7�������w�n�T�׮���s��I�ܱ+<��عE;޹%�P ���(G�j䀤u�; �o��?w*�j�Cȳ� �E��FD\85�7(+hb���U����N�6pa���Uq�O�ߊ��	E�:_��z�V�i��m���>�(/r,������o�Q
�Ae��*pJ9`�y�tq��,��bo�X�vw$4��>��l��Vޭwn�~�H�K��`}�N۹����.��ll�=}ԏE��_�o�O/�{�aBPn�)[�3�������UIE Y�(�	��/�4
2�˻6�qˡ��˫o����x$�%�'Xz,�33��[�eT�:A�)���J�(D'7gC�u��!Q�)��yMoH=!�D�'����L@y�9�h�����=�����e1�2a܎q��a�l�Y6Y�qK]����+��N��~��]p�iz(tV��3�*ڸU�3�(�eA�/x)g=a�T���ԏ�g��x�]"^��qxb���280n�)ư�c��j��s��k�*蒲�eK��yr^�4&r��?~>ܻ�XFս��O�n�ٔ������?�7��ٰw?<�Φd=0�u���PƳ��y~��i,��B`?�T.���|��6:"M�x�_	ѡ�3O�MOt��-\n���훛�����5���T�����<�舉�>K�����d��9}l8s��p��Q;wb8t��� .*{?��\��L2������1�r��&�^i|�����)�|��/xO�m�ɇ����>�O�֤Oͬ$Ԅ���s���C<^�d��p���޽φ��N�ʈ���.^ĸ�E����% ����qL�q��8���fcz�j�"����D�?�#���n�w��Ƚ�������!�Վ�o����z9�nh.
O�8�w���} #��LŸ��H�3��¦�-z>���M�^!Yu�����>c������+
���^��v㓾�8�G�����b���>���?��f�S�gz�(�<�A���"�侟�����.4�~���S�;e}�+@"�e��f�3' �HMO=1��.@��=�h��>�4�jJ.��P��]������~=�����.����8�#�Rh_�7�� ��3�e��E��
���!~��V`�<��w�Q����T?_G1bl��8�G/���0��P\x{�S^����RV�N���_~�N�7��4:�\'w<�_{,�F}�7n�΋��"���uu(�k�������1:d�X�:�A*>�4�ٸ�q[��b܊�x�.��x������tdF�B�Y��MDR���V�HN�OB\g�>�q��5w��i�x���î���_�����_
�PB�����,�g�`wT#�g��̭&4(���ؠ
Eс�.4|��!U��|kN�aئa�E�-F��������[�/!���')^���,�g ���#���p5�eZ6�ۜu���
q��Hr�oUAL�ݠkn��w~GF'��R�Ը%Ė;2u06~�� �:)uX~:���;$�yV�؎	M��Q�ˏ����ތ�2���D��ܬO�z=�:��7�-y^�E�!ǘO��ۥ�F�����h_��=�	ࠌ/^�ş���7�K��ژøUv�R��Ԅd$Ef�^tda�K�=��A?�5L��7�x��6�B֏���l>R��s�A>{�Pr�U�a�O��?x�Om&�0n)_��`��JĄ�7���5h˸�*�Q
�@�\�[o�>�-����3�����ML� 	�K��K��1Rz.�g����7llN�>��S|�yx�1t:��������wB���{�.�%��1���1����2|��=ڃ�\c�#\�?}ΫΈS&Tb�#BZ�U-+f��Ϟn���P���ر��Y�W�\��x�������L�ַ�۸�s�K�e�mr�Sw��<�m;���������6�0lٙ��fA��_�x֣N��[�k>D�g8{�����2D��/_ø展�����G1��NIyO꯱��q��1�����>�	}�k���/t���_�_���-\x�[�1�u��J��Ϟ<���xux������-�9�������?u�Q�$*]�4/yc\�����(^GF��[�M!a�Z��֣L7n�~��/����_}꾷w�!��'Z�/zd�oi\drS���b�׏�u4��0L�~�8��,gh�q�[E�l��(B��Ep4�16,����^�uu+]5P�wn�V��i�{�S�O�h;˟�nah�r��|�ӈ?�q�u���<;���h<HJfכ8������o{����dt�7������2\7dd|3NrR|4_�k�;�6n��pܹj<R:k��#�E<��(ʶ$.�O�*'�[��z΁
"�/��K���gZ��k�x��n�p�̱ᝫ�]�������̗���EYb'1'�ӏM��d��$��Ү҈L�F~��Ê��(�H��F-�xu��+E��L+�F�J��d���g�:��rY6�%
7`4�٪��!Au�\�i���ӅM�;&L*�MV�#��<��I �HC�%�L�,M%9�,�g�#��u���6*G���L6�"\5��x�rԳ7A4/G��ū���ueƼ�=~Ш�e�Sƀy�P�\%�^�M:=L��xj%}\i���<�B�(����!zV:��;�rG�w�F]���"m
�Y�X)��-�ջ�L"��/�������]r��a4����ӄ�Ū����G2����Z���#[M�Q�(Ç���1B������^`�2�`�<�M�#��?߸[���Ɵ��31+�:�����86�`�2�Ő-R6�(	ԅ�ZH�"�Y_�y�Nj��=�}�s1=4�CѰ��arƈg�:r�r��A�D���Z.�:un��'s�9�� cJ-Ƣ���n���`�� ��O�����E��r�K�X�>�����G'x�U��d���';�b������ꢓ��'8$��%n*;;-�ԇi^]v�ޣᮌ\>��g��lJ�1��`Y4�\��pX��NN��5k~��/.hg�]9�d��Ԙ@nE�B�'6��ܦ�a�G:��d���\��?��v������-��e�m-f�:
=Y3>�C���)�h��^��H����L�D� 3��?��+k��i�d]b�E��&�A0\�Hv�Y�QO	�=�ڧ��q��p��餿��C��`��<
�O�j�ڶQ"F"�EֹqYlx�.
��w\ek�ۤX1l�c�y�m�yN`D����/�ώ�'�h�ҏø�<�'�A��D]���<�s�r�.9�I6l]�UM�G;0�Ņz�<�ql�wn߾|��[	�KW�,��JQp������d���r��T�wI1 �O�(\D락��їR�]Voхq��i�h@�
�+,>lm�5`���'���+�,��EH9p��[�a��	��JSij�Pv;����Qn!�x�ڤ��'���H��'�fug`Fk�Γ�M�F#�D�� DZ޾��7����	P�z�g�0r�[�:NsM�J��	3U>�V�x�j�Ae�ǻ@r'��63bE��A��0xya:�Y��"�WҺ?�Βˇ��@�0.��4A�<��;D���_��f���##i&�''v�t��?p��g䰑D{��6�u�_)#��2]�wT͍�^M�*��g���kP�I#�[��1�>� Ѯ�
8�w��Ӯ1�L����R�ѨU3�3� Q-�d��0�h3��)�6c~s<}�ldL�AƩ\tk���m�+u�1k&�K�B�⺊Jvyr��2f�/mlj=`��Me!�!'��sE��k��H��:7b�}��Zk}��y�Kk�(D��b���ݿ\7�\Hq�/v�(é��hɏ#�	��#�v@'(ϔ�;�5a_���Gm���E�c^w��{��͐K?��V�*��%y����l��9X�9�3�����.<��}���s
U��?�i��^s�b=���C#��	�H�����%�,EgZ,^��%�_R���/L�6�}�����+j���"]L=���m�r��v[���7��ΙX<cc���b��W%j��q�t�Gv����ܲ5�Y�!jb�и���Q�y����m��Y�'Tf3n�82��8G6�D]�v��q��3ǆ�.�v�g��������)���*�y	н>��s��N��4 �H��PQ1�Z�V��G�u�2��q��n���-�Z�[~�a��-��,���C�J�۵�k!�!C��c5yjaf��	v�����Mpgg�l9�(kX&9�8��Y���ːLK�^���&���8
D��؞�d�ч\�<͘��)�&�L�H3� v\|��	0���|-N�S�9��`"A�� �Տl����<�L�k�.B)�[��l$p7Bc4�y#���%�w�l�'f=�ayYX��;\�"��%��3�s)��+�|-3��
�c���&�S�4�`%b\���'~�����k�ȋ'#BV����F|�?d����,�8�	"����e�a��#(�,�����:py�sh-@��*�;�E���UH��S�YЋ���1E ���B��8����U���rٲw�:���:sQ:ABӻnr[��-9�q��h"R��L3y��ī�Ug�JS�9ʌ�8�)�dG���}��k5}-uk��@�B,�6.�:�|<Q��r|��&M��]ІU��p��°_S6`I��%����89��wqg�heV�-=#PH�鋷��C�v�24}!GdJ�b�Mfx\���^p���µ�'�q�K�z��g�<+ˣ`{���^ޣ~�wVO�[x�y}�ʚ����/�y�6�[�>�d���K$ә��6n��Y�.(m�"��6�m�񪦢��a�>~�@���ؑ}2n��q�?�_�_^��h��U�b�Ai�S=]�ԸE�D^Ÿ���J*�V�z�
�=(�|^߸e�Wɵ�q+��Wj2�g$��.�t#n�Z���CVw�c��a6S^�ɖ!�by��*f�W�Y�c�򖑅���"��-_!�fLț�%��-�3����O-FE��~���C�Z\ح<i�/ŀe�� 'gf��2��y�G"c�����(��c�4Q$"d��r��a	?��y�NQ6&Ex*�\i��P2%d"����z���o��c^��qK�՞��d�ב� �5�W~�G.^Cy*�`"�J��	-�
���Yo��|hT9���.��SR������]9��Ӗ ������R�U ?L�%
e���b �,<ԉd[�rڸ�1�Lk����׃y�z(�E������c��)����9�z����E�t�r�x��y_�㱘k�
���Vc�U:���x��qGyB��E�΋�t�$3�6$�.��gt���Vz��뿠�k�����5���������G��۾ �B��g$
��yF
� z�;��!�u.9�K1���kt�3���uƭ�'�b'��Ŷ�^c������6n`��q�z�g͸�>l*��~��5y,����E�V�(=���()��bc�8#ko��Yآn�`=3n1�øݳ��p�����#~,A:R%E��`'�J�����?�spˇ�M��b �:,�:����J��Փ),�9W�������.��q+ �te,�����kC�Q;j�gQ#���J�q�IɃ5]�T{��H��G�c|��r5�{?iR�wp �dФ�d�չoE�b�>��܊�[��w]��y(��k�u�U<�l�+Z�8��v�f�/���8��}�&Ôߥ���C{eZ�W����6H�=�NH�i�VP�t�E��hW�U��}iԳ�Zf!u��'�뵀J�\��ȶ��G|���E��!o�(S��P�xd,ћ��E�ߖp������%�w x�΅_� K����d�6�>���?~i��H��S�лZ��Ȯ�p��V�uhn�x�����Aخ���E.�����6bܸPn*��
A�?8,�:9��e��1���
� 7P'a���-:���B��t�;!g�S\�2e\w�:�`�K���ƪ~D�.���q:K�ɹə~���/ȁ��3s�
K��T��?�+�T���cB�t3��[�#��
]F����V���at�J\,}�#��{�n[�V���+��0lF�vK�H�F^�Zc@������V�"Y/M���9��%�dT�g�8Ǝ�4bˠ+;:g���^4�7��n!����,����.+ഹ� �{�����T�S\�7�zM�����$��.>�/BK�v���H4��%��0��S���U$����O�,|&t,�Qـa���3����0�V��4��w�iୠ�2bf���,�k�q�)(��n�!:�E���vp[�좉r�(��2�(�4�U��G>�tX�Am�]�����?h�-�G���T@��W���a�4�O��m�����w�q��������[���zD��J���5 ��T45�e
J�����^�v^/m���c�Q�q0%��eH}Z�������mP��s|��\�
J�Wi����N䊊�
y4YF�I����vy�i1l=�;be[_P%�4�����;V��l\��\\,��Ā�+Ɛs|VR�|�8h�S�3���<\m���8������/���������W|��(�m���gd���qgGkhgU������a��DO�F����^��y�<�Yv�N3Z�,L�ϲ(��=Z��L#��E��Y(�5:��LO�8}~N����Sh��R>i��c��t�8ʲ���D/s~���[ԟ8���*�2�1f�\�����	o��|���:꬐:bز���a����L�X�(�|�[�!Q���i���(��cvQ�
�A猢5���0�ycO��l�����p�?jAv�}�!Ǖ�N����֙d�
������=�	�]�Tq��2z��u����FS���[:n�G���*1�}@�*{[0���R�����	L�Z ���RB7+j[H��qzy�]5T�:���7m�ul*���˘�$e�lYٵ���%0q`�o�����Q��<�9-�:��$�)����`���eM-��x�����Z�	��	]���*��ΉgR	��S�+��;q�Z��x�/�k��\(�	 ��<�k2��-��-_�H27z3G�Ϫ{c� �SG�h�&88��¤���ۀ8��vh�w���@�@�0SñW�pLy���:�4�s�H�̫P9�Dq������[�͑��~;�w>��`�N�h����S���Q��Cl�� �@��Ӫj������Tt�24kǵ�o�YF���S��0qI[E�|*��ef?�;O��gZ�B$��*�c���ƾ�R�Wr�qܮ��V�:����`�4��>Ê�y^�U0AOI!UA<c���+z��hӍ�BSt�6�cT5ȼ�s���f��[�]���3�v4a����l	!��"$��˞�����>�.=�łʄ��ҭ�)W> ��RL'��'W�
4��够��"{�DY
C�!�0xd\�{' �̃mhLF&�x��J�I
?��O3�r,G�0/�+�X6~�0�,�'�<BtȄjȸɊ|�s�#3�^�Y֠N�p2(��͈��]��IH�k0�*3��u����58O�������}��<�@�y��)��ג�:��ś���-MR��M�����e.t]�q�d���*!�<�j㴓�B�=@����A��@�K9�S"<�Ɋ� ��AzЄ��F�q�)T���Z��g�0q��c�9��a����˗i�߀�fe]ဠ��y��<S�帋r�Ү�"�o�u �>�$�(O�\z�V��g"w~��̷����k}e�~.`t3�7�x���w���AN!y�OG=��1��������E c�q���uQ�O<u� ��#�1W����9��N�+�9r���>s���B�3q���7'D�+�*n��EX�I���8">�*������˰.=[��9�QgE	��Ǽ��^��_vǄ���V�1?G���o$�Za�����#L.������/}S+�_�mx�R	ﻓ����q�������l�2�7ݔ�<�^*�sG�'����]��ܬǢU���<W��;�82��_���Q�c��(���Rl�\��@L�+�\s�Y�@��qG^�Ӳ�%��m^T@d�Y����>���O��#F糧�W���\�=Ӷ�<��m`��A��g��������I�gX����y n�\\T�~c[6 MN�����~�d�֧ׁX�\�,ǻO 2W�=��"79t��2���]\�U�){pN��:��Չ_��6�"�M���p�N���uPI�O�ak}$���X����\\Z�w)�V��U9Ǝ��uS�`�I���5�s,Js=;��ѧ#yD�ci=��G�wHyY���r��G�J����)`�B�(G�
��X8�NsZ���r��F~��ůa,��u
���E�A:5Dy�� h~ e�5���fF@)S�V�4�ʓ�
{��dI�瑟B�SW�I�2Ƕ`�)oQ&i�PQ2I�r�oUyz:CK�J9M�Q6��@�M2���Q<��䨚��N����)�a9#�QΫA�7(k�M�;*Ŀ�s@w��p}=� �BTJ�+��J�f`9RI����g,1ư�����}�*��#D�5��PyS'K���@���(�aTP�
w
[��Ê����V?�	���<W��1�$F��pE/�j����7b<���q$�W�m\��
Ð^NKd�KCet��e����ZI�3�#���6ް���1m�_C�ww��&�h��`u|���Б/��\�@�g�$<G`)�P�ԧz�~��		�y�>��7��q��:��B�]ۮ@�����D��#Uϳ�Xϳz�qPeU�&^�#�Ф�Ο����:t��03�)������u]�A�f�_�m2�0i��a(}W�@8=�jK��Y1�L�
�#X*���X�#P=j�5�K�Ú&�Xc5Kr�M9������ �-��X��cuJ��"LdL�9�M��`���Ce'v�{�X���2�/�Pe��`g���b(h%�P�JJO!	���6�j~��ؕ�:{!#�;�[��|e,�#�qE���A��w�>�`N��&�h�fy��Nk�Oy�~ �A����[�T˯��	�V\��#�`[�f}i��e6h̃�[��1l��*��Z�����%:n=pSw�О�|կ���U�������4�ə:gi\Y�;}��2�mL��H�i\��Qw��t�2HzU+�4���^C�����&�X�Jr7}M�b�-'幟'.����kҕey�\ѷ���6>�o�����	���k�x}�o�ĵ�G��]	n	T�'� �\�"��+p��4嬍�O��ib����X��m��5�DF\+W��2��O=n/��m]����	�4L��ݍ՝�|s�ۨ2��[zk��-\m�%�;Q%�3���v�u����ʑ_Q�f^���G`�8���3�Z�%W�M�NS���1��)�� z��2	,`�R�<�K�H$����B`)�G����Uκ�֟�5�S4���<k0�1��b�;	��>�CO%�IVc��#q$0G���[��ᡢ�����n�<�dx�l�?�,�a��ی`�`�K?CI��E����<L� @�j(��M��ǭ��8mDe���mH�\V'y� gF}kྙ�E�"D�؄\�hpz�"c�)��"�eKw��I��ʁ���<o[+
��ޟ(�(��(�S�"犘%T�j�+�T9ۂ�qZ���M��zc�zXƉڿX*�0��d��?�7OEt8��r��Å��2�p��#o��Gچ�2�M�icx�g���a��k~y&|*�r��.�+_�t�t���'b{X$k��8z�ۮ��t���ߖ�TWK8��B��Ú�`>��cY7��ָB���ӄ��ĘF� ��ʯ����.�tx����{( VQ����/o�Xqrm']��wN���;J� �H�z�?�+��T]���a��^k`:M�q���΅@�7���ehm'�UxB��;jˤ�q�`�-�ly$/�`��l.�}̙~' d�
t��BY��)�
Yi_���� |��E���q�:�(:2�i6���Z^Ѱk�l��D����
��r���:ѱ4q�Pro/?,ɿ�c����:n�@�s(�v(�٤�{XWH�}x;���ۉ�.O���hۻd}(^��&:$��.��
ێL�|y����/E-^NM?�FL�4x��lD����$�KЧ��)�t��A ��S)3�i��,��a�D�ܪ�Ȁ�h�+i$th�鶀y���OL@4޵�줖qW}k�_n�W��'�|'�Z/����W�-q��:P/c�Q����X��kbY�b{�D���{�����Wh$��&C�� wV���|+��U7��z��kqw�����р[X0��U��˘��+5����]i0�F��g}2�k�&L�c�8�͚5F��Ҳ�8�'}�����<k!�,��׺U7��am��*�tܘ����/�����Ѽa��[���JG�'(��nbA�?:G��{�BE�ː��g�I�7~�d���2��"�F�������Y��З�ac�+o����Lc8:8���+�:z�vs�2_�g��IdYE;#�z�:���Iڴ���@�;XC"���4.ꑁ%����N������ںc2�M�& �A_�1d*�J�E�
ŷxO�c{�:jQTp��Nhn�{PT$�g��������*��+,����4}�R��#4�>�� Z�B�q!��nmm���'(:_�M��1� �|S����RTLk�_�ӅS'+�b�SAɽ�bsT|��Y��,���>��%W�%t�k��E�V��kL���d6��d;)@�{��������A�����ɤ?`X��4���ep�H�L�.>��[g �QvW~��$��r�<����j���1xu��EA��타���N�tz�/��m�a
�}ԥ��ҁ~��!~���=>�vT���:�̖P����D��l��s
z�nʇ9�h��`I-g�؇����~�/���C��ᖇ����h$7B�c)�W�2�y~���δ�E^q�E��1G�	ZL���5�&��W��#�Q)��r�z����~�C%E�+��"LթQ��y*�#�*��v�Z^�yb�N@E �淮��s9슶�R��Ǻ�S�$_c�V�3�8��"ɾXhwGeu#�m�>��bA�Y�*jLK7a�ZF�H�ג��#��P�U��S҆�'f�@�Wg!�J�]q#��-���j:�.����$	��#��V������<�I�3 �h��EL�2���m��&�}��Ȃ\��S~�j���s��L���.���v�q-�h�U~�+O��d�3 ]G`lȕ��kq�Q�D�4��7R�NrA8��8�ve���7����H��_q�p���j��X�V�+�S��K�4�9��������QE� ��.��:
�79X_&�Ե����{П�7��x��YB���-J�	���^�����R��ߔ͝��Шtj:�5q�;��gX�-�Ec��!�D�s��&�g�`�@~ʱO$����]���~*���f�^�!y!�,#�qt��a|��]��W����##����ѧ�O��O��E.���ܶ�,�r���~3ϓGz��h���	+b~dB>ezIF�A����DU�s�B���=�D��5���Ù��Z!3s����>Q������ٷ���'Hu���3��2:N��T�,a�䁿\%p��~-�!hL4�в �ɟ�;��2��<p#��#c`4�
��!'��R�Ϟ�*c�S�BA�^�oLM�Q��r*s˘�(i=��Y�3hzO�:-C�di8�E����P����1�N}��?Ɨ^�2�e8H8H��v�k����� �xc����W�Eh=�đ��J�����y+_�q#J(����:.��5^��X�ʜ�y#�RA+3��v�<?�_OR5̣꼀JN�S����qN0�k�[��l�lq���X*�~*^Aԓq�^JVO�Қ�.�製?�C ]�~ć �T/X�6kʲ<��^E� p
9�%���s��F8��� ���i$�@Ҏ��$뀒=�nGAb �-l�6���.t
:y��R�ٟWq��� �-�-R���h.85� P�xb�� q�P��G���\�����o�,��9$����1M��0�e#o2����nr�Y�[\��X�a@'�E�k`�d��
 t�+�F�C�j�D>z�E��r"e��gY`}�rAE8�֕F�!����%(�F��I����#�Q~�����P_C�GB$�_z��\�\v��ќ�'`R�M��Q�]ad+n%�e�nU�]�W�W���!���Ч-�o��}P��e�7�ψ^��Qē.��f}����*�e0$dZ�.�ĸ�� d$>�º���F��lE:���Bln;�	������ ��6r}�ǪO�@E���5�~�,�����B��&CH�m"��:�vJ�Å�g O��<V�˲�;��D?�S�y�!"9��ZV@YK's,X�ז�F�`?c������è�:hP�$�����_�q���_h��'�iDKP�ь�*t����aZ6������	���-�:м�9u1��1�q�l���P?�J5�xd���K.(ʩ���*��$a08����(��c%.���@�cK(�o���YAN��
��Q�j����:e`
f%l�)����o��S�e�eY����XC��1�%,w�Э����@ֽ��&3&��T�5`ө��	vqQd�nU��Rߛ�m�S�
Z�q0ܦϮ��Q�\�
��� z�@��H���-�j��i'[���SV����.�$q��j��C�w��'� I_��������/v/d�>{�L(�6�ۘ+E"�Ѩ��\�I�'��I�v���}���w*�����d��x�P��!�_�?w达-��]�t��$ư]�̑���	g�1Ih��1#-�/��)�sM�E�`[�"X�![@�^?��U�&���fa��D�k�����9�~+7Ù3�����zTo���^�+~>K�7?U4��Rf�(`��=	��ׄ*>�nW�밯_"��]���ʀ�綛��ФP|�K�xΫ���+���z�F;T��B�eg����˞~	k^�* )סi:\I_�)��Y�����:�"�[a��5VA�ժ��U��c�!���@�F�uб�p�<9Y�ĬsF��"qμ�3pt��Tq��H��r�~��D���$� lʿ��'P%��ń�e�b�E����n�d\Oە�3���}��-�@�3�s���Pa��gO_O�<b�ʰ���i�|�o�:��l�ޟqC�F��L�ؤ.;���A���q{p�`�,JOk�u����x��6���.n�:89N��A�.����ۃja�G`�V�Hc\p�WooP�S����)aH�dȀ˔�T'Y����cg��M�P���UZ��ZPeX�%K��?E�Y�������-B�a�Mg�Լ�@@�NF��~����!�@1��lMS�%!E��+rOÎ37C��Ns�i�W�(*p+p�Hd99�r���4��Pת�R�+})��,z}��! v�ڮ�rPݘw�����7KU���`K1��Pu2��:f*�  ��IDAT=+6|� U�0��-��E�5�ʝ�V�gI��#���+���6^�;��{�y����4������n}���!���͋��g��ڰ��[�s��`�����mԦ�[���6Z��8�7��x#�P�qT�۬`g�e�(S�c#G��	W7u�s�)�:*�-�W��Wi[� iH~�z�{����3���.�4ݖz�f��7,T R~�PJ�bBKe����T�{%pU�u���o=[�2���)7
6���c�O@P�U�$}F�z F�c����S�lԮ�1!�2cL�qB�:X���&�Ճ����a�d=\K���4�D�����)��[�'�)�$����'P�N/0z�'����uv�y}�A��w)GÐn[p�V�aֱ��{S�d���c8i֠�n�z�v�Ώu��������4�:�B����J�\�{.���⑄��49�����Qa�j�����zP�k駪�	���1�d=}(�b7]��8N�u��Ҡ�7>=����yiQ=�}q�Ȼ��9D���͍��ܖnUK� �^$*6t��S�����*��b��������W��mT/!�3�P��c5T�����e��P^����t�P�#V�n"�0~��r������
C!����\rɐT{V;�����t�⠵K8㖠�A.�&��A�f�rv
M��>`&p���������˾���Y�[���y ['��vR��v`"���E��AYFr�	���2|SX)���6�K=YW`��Ip~_���R��@�q(���j�Qn�E`G�* �-�7_S.c���c���K�ڡ�9Sa���9����߻=���x*�~֖�S*އ�G�E��;��E��JN�&�������� I����"eGus8hO��G�-�-��d����m�&��M������ @翪�i�S~��T���3u͆�� �\��댯����u�!S/W�5��(�����oK�cX�7B[�D娍7��P�c	$�h���7h)�]��^Hh�nHa|&�S�Oa�|
.7�/!�AL1A 悜�m���yu�s.�d�DZ�\e��mRHӁ�	�=�*��˻�Y��[^e������X�d�#�� �$Qy���G�F=C�w�u`:��x��--G�	i��h�HM:T�M��Z��s�`:^��
�\f��K���Z-��R�.������r��2�`��������o�ئ���v	f�_`�.ʈ���c�<?d\�Ӈ�n�W�{�*��2l�_�)���o9\'ƄЄ"M�"���{TG]j��@���#hZ9kpK�|�'��!k<Tf��ߋi��0����-�-�LU;�k�>�G��pV�`n
]�|F��l&*K��$N��]���s1.P2�Z��V">�'�2���!iH%��;�sK(V#�(5�U��L�j���&�*�Ap\��:ȭ:�:�:�T?�:��|B��)8�E)~:�	���cA���]�"y`��<�����(#l��/�#��=e�hՓ|���o�vd^�-S����"�3}�:u~�U��u��9E���0ֽ�d�3F�<�9	z&]��bȂ�+�:a]*1v��):_˻`��l���.��K�F9G{� �*�������S�;Q '5�;�:�0HF�߇��9�pF_��"W�s�b ��9�OV�$�'&+2a�+�t���D�iZ&!���V�GY��}y+b� "?�%vǬ�W�!}oB��-Xh�B�=��cݧ�T8�T���X�Kq�	��j��RX23�5��TZ6�8j�o���žwUn`���X��"8Qo�i�f6�~c2b3���r�.]'������!
�c$Ht��:�t���&��v�T\��4��m	N��C�o|�\.eu�c��۩\c5g��5���o-c��8�՚Lz�K�&����$~�J�j�P�rY��%F@�f,e��":E1Қ���o }�;މ?�B;鮁Q�t�XG���}K��:�Ey�Oe��wSho Z�-���A�8Y�����_*��s��2"�ܬ*U�r����p�	�M M �(>�����O�v$�3l�s�rJ7.'�����^��#a������+��cd�v������1��7�Q�W�7����3x%y�0/b�̠$�$���Z� �=��d�:D�����[�&�Q(��c�N��,U���(p}{������)��@��9�=A�m�V��K���"r��rͰ�z�Ǟ����8c@�wD���{���� �)��BG��"*��;��l��>Ǹ�lׁ�Y�#�0R6�P���hdL�
E?��>Jk}ɩ��8��0�,[ƭ��.��`�,��hDaN:)���"@u�v��]n�<������ϡ������*�gk0�:9����0���+�ȩ�m�����{᭓iw��W�k�T�W�ߦ���*܏��W��N]z�>���o�
L���.4���o��Rׂ<I��:A��2����,%��v�Mm�P��N�R�,-�k/�)�U��SE[欳�tV�W�*+[�i��-��W��ts��� s?�7b�3Py.[�����6l}܍��|��H.�E0�(��k��Дa�>���W��B��!�ʬ'�1z�= �^���J�U�NWV�u2�b}�B`�Pֲ�z����<�12X �I�9�<y�GD����O%�9Ӫ�: �')5�mU��9�R|�d�j!}����M�YE�nR>'��5��S�ׂd�����2�"����Pslk�T�֦���9���ҋ6�l��C��^���;�d�[��a;���\���Hy�g��3���������=-�.�N�wچ�.��'�T���|��aɧ��U.�[aO�y8��]�ج"z���H��uՙ5)��os�Ή���[��fNҋ�����0y]���!�z�m�l�?�B�}��r��1��1���� ҋfP�(�> f9f��w
!�z�N��^Se�������%����n�p[�����w�Y�9�Hc�C �2!yFz��{��&AҬeU�0l�� w^w�5�K��q1Y�W�ND�.���*PE���(�V`�Û��U[�l�B`).����Ǐ������xAË[��������@�y�.���I��kdئ�&w�K�=l÷�:���#P.�ǫ�tw
5G�oH|��s�W��0�F,�D�p��x�'.=�C��u�\Gc�Q'�1Rn�:m���w'�y�/f�Х�G�A�1������ZyUVb+�ҊKô�z�.���z�����E�z���:��z�P���r]g��_��-���^�1��P�򭢓�1�?��4�'�CE*$u��mU��.�W�y��K>�V���� ��ݕ�vpJ;��Rm�G���;�
���V�z�\ {.���e���-��v �+AUu-*�{�ul�)A��Y����;�V��۹s�.(�� �Zm�^��������ϔ%<�5��㊮p�S��FI6��"���'B�"�|�W�R���m; ��:�^�dw��z�e,=��R`�0���$nd��������7�~#���B�js���vm�Ad�ǅ��x�>���� L|�G@�e��5���<��w�%�v��a�F��i�4�,NO�<~c0�U�UV�]Bi�Gɚ����m=d�~��l���7�@EJ��-�<���-՞d&�ô8n�i��;�̷�s��䟪WBV��Gz��u��Yױ����8�PU�6�� ˻��rk�����<���*�C���a	([N�w�e=s��vG f��V���;%�s�N�Z��	c�������k@K��s�L���U|	8�rVT���P��db0m#� Y���',�N��<��I��K� :��ϊ::9�2"��X��MqF�`������"b����&��6A���{T^�4K�����ʬEd!v�:��ٍ���x�����w�3����AO:�Q:�p��@� D͡��X�V�Ԗ�rv�8�'��dL'��v������)IK0�FY#m��H[�4�ZH��"_K�ӝ+��},Ɩ1��a��<p��FSH9����>�[��4�W,�%�̌��g��A��-��������J��YN�3G�IP��k��o�_��(S�W2�i��B���|����Yqk���=
�u�%���]�B{��+(����8�	Ζ���2�v�b]M�W 1�G�-n�G>^�6�kQ�Iw}~�� P��)�.�����-�*�x���GH^.�����/@W.+��D��@���}{�q4�dc�� �o��^B'吗� ����2'�NIb���RmWv�J�Q���:�KR�.)�	". ��1����!,�d�bC���e�b3�òS����������Trz##����'��?������9��
got�\\B@�8z擂���3"D�\�睎~����<1���/WL�U�~L��u��sU�xِ3���%��F�fLw�Hyyf�o���~��ur�#�$�R��R���hУ���a�4~6l����o�ɯ�qT0YN�L��?s���ob�+�
")鍑f?M�� }�Y���5g\��Tn�$�c�ZY�i���F�Q.O1��#�f��uDT*CU��W�wG��@�J�#
�O1�
M�ut�(�x�t�w��$����2�C<�]���_�.-�	"�)濉�>p�wyV��?���f���*�o�����3�1B�A�A�\�Q�༸�+�g�8p�W�SfE�LGKEc]�$WB`���I\
�o8v�
�5O��Uӗ��뱤yL�<֩�ɩL�u��w�dp��ƌ|���G8�nɉ�h�g�u�Y��PH��c�!�E����Mw���',\�4$��h'���3�?h�8�p��a�c&cO��p��9�\�b{���Ι�L�Q� �̓p�I�N��Dۡww4�O��/y�Uؼ"��c�Q��4�����\�M��^2��H#?\8̏�'A���я��"���<'��$��dx�H�@���g����o����AF���>M��k� |Xc���n���e�ʷ{�x�яǓ\�c;�u��e[�y�G�}{�ف������i�4�,>ϟ>�}�<�ɺA�<ٯ�+������: �ʑW����ȡ���L�7$MC��
@��VF�@�.%�G&���)���Nލ��І�WyU�ą3f�o"Ɏς�������G��� �݃X<�o�C�Á"pV�%f��`��l�0p��§8� %� ��bN|�	�m��	'g��y,cId���*�r��
����Dخ��W�9��C�:�Թk XL���ē����=V���6b����ÃP���R~�^zp}�V��g�%=y�������v$�Q�D�.l�=��:��
��=���?�0�J�����AS�Z�����,j��+®��PyS7����H,�9Pp�>��J�萅�8��@��<s��d��k=$:3�50O�lSP	�G�*�[?f�]��W�ҵ�F}y�
�D�A�ua�߷g��S�-y���oIᄶ�#.����� ��M"�� �n
��5^F��8ו3a��+�4F�7�����i}��g�t���\8�wx�s�B�x��J-�LϨ�D����I���%o�~��h
{Pl[�3�DP&��:���w����i~9�q˵�HT�v�_u�K��.r��l���dh����5A|@I#��H��#,@�U\�ў�]ur��#h�SP�۴A2sF�t4��:K���]�̠/׀�:�
7��*۔ӫ%��z�B+�q�Ph"a�HI3���Z�xu���������m���L��+N �D��h}ZnKo�W�N�S~amف���,�ɕa�v��EI��t^E{w�+X�s���}���v��,�o��j����P�+���ǵ���U��?ǂHi�!,���5X�}��9je���"
��X�j�5ĸM˩�<�/x��A\�)��8m	�^�Kax���-���Q�:�wYF!&��^V �P���[AN}��1�:��q��ۆ�"�c}�� �h=�����C�SȲa�f�|WewX��%bɵ���s�P�˰z»5�K�s���;���m�V?q��]s�� ����g!�N��,����<㈼Uz� ���|:yLT���3-��r��t���;��[�^��b|(��������;�ɘ�0ҵ�� �¶���|be�]���
u2F�
r0�0t���8��`!* �0\c�(y�:Z��$�+�r��1��N�=���)�`�.-^���#�Q&��N; ӆ�;�m�-�u�;ŷ��v=�
/�7��6-�)��aZ��t�>���c6w��}�]Oa�~��e�<�-H�8d���;_ 8�@+��B����YNe�md�e(�2��*�s����c-����w�H�����(�/v�V9�d��X-
&I;�� K��0������i}��^�$F�׋9���_��:��e̪�^�����S\ӥ���c��k������.��א�inٸU������+�1k��Ǝ@
�X�;f�spS���+o��]���2r�0�4[@ucƩ�&�낸d}TG�(�Y5\5�o���U���8�O�$�|�˷
�
LhD�1�dv���5��-f�f6�1m����
�㶰�I�<��J���	G��.�y\�=��&b.�<���u*�>���Tz����;@�6�.3��h��l~���2H�y����20^%M�3��o[�PO��j2�L�`ܦ�^�U�/�S�v	uJ�����P���栚�n�,��ʁ�TG|�8O���բ2S누ӻ,	�żpYL[�mW=�#�����0�N����s\��ыm;�!:G܁��aس������������:���/eܒ�<���g�@��;�M�4��e-����
&�Z0��E�Q��d|P�y��p�ϔ���q6f�_�FE��@���n
GT��2T���I�K��0jK�L-�O�}�R|��.Vr�4��;�����`7O��B�Z0ڲ�B��4^���-ibJ�Z��ذ�d�0� (ل�k��-��FE5�ZR��t4�ia�$��(^sLW����j+�ʚ�Nr�:t��}�sqVͤF�S�`�<lX�\��0=)�(_`gL���:�>�&_�:.U�?��[GY���+�W�Y�̦={�{�	�7n�^���)
&EW����� �A�� 빨�AG�v�9d��T#��_Dj2,]m	��&��P%�r���w��-�=�^Flo����S0K��q���G��h�	���m��K(;A]����Ҟ?W���͘u�sA�7{�W��.p*����.�+f�&{q�#��S����Lتg�������ο��tJ���=�Ø�y�gȈ�����0u�m��#XA�!1"���ytN�C��5GQ0֟k��c�bd�� ���c
�J�3�"ltٽ��F <���B�@�*�X��4�_�1���� K�`)��.��`4�f�A�S�7n�'_�[%0�j�g�@�c��۷��߱ �aP�e`�
f��9����
�,�с�e�*����t�wj���-�Y��%���k�3����Z��,_B���ʥ<�?&q��.��ުC|������&ۤ�Ul0�w�������tׅ+���"\1J��\թaKK�Qj,?E�Tu�pϣ�,�E�u�X�.Β��P;����fj;�/��B�&n�7�l�R��fyG���|�f�V�n*C�q������d/Yg���L+3�V�I��A��'��˻��2
�_����c�iAϯ?�6'6t�zp����t�yd���ksn�W�$fy��e��|�u�؂��PX�˰N��L��D��a�F^@K�		��5��|}������+2&yp�<�P�Wy5�B�ZZ��=1y�VPu��X�@�OOp�N3���sYD�
|��W�X�[=������H��.q��Y���C�6I���
#Yg���5��@r���p寴i�������N��2����h�ҙ����\��r����n������أ��[G	��OEط���a���U��DfS��(#��!���p�n�oq:�>��ͣ�v!a���#
�2qB�Z]�a��� 
�~�i�,�H��ir3>����U���]�)��y,�a�4�|\�?�]¾����G�����[
���}��V�M��%�Ƣ �D�#�8�+/I�����u���Qqqh�2�p]V�����~Oe�b�OL(_��c���Q�uF*N�H�CWr*Zu������f���u�r����(N��/?���Q�(G��Y��`
g^�%��-�K�LMgY��/��j:��t�O_�1�;\yL��8�8�4D������@�	#���q񪾁���7��,}|�:-�+\@��pjѧ5�y�d�5��a���H�'����-��1������-��RwS�r��,����}�����ٳ��n���e抮�9��ͶY�/j<�#�M�GZ�� ��逮�O]:̺�P���u�����/�N�:�Qƴ~=�s\�����&��nB?��BǬ{�^*D�`������mѷ�m�3lb�α@��S�K�['��ve�d�ut��	{�I�EǑ4-��E)?�{��������o��ͨ�(;y&D<4A?BŁ�V�X�A����A�.�q��i��&`�v���Á��e�ʸ��!�(��D'#N@Tt��|��y����� 2� k����e0���gGR��}���.�7�i��PyS�.;��0��S�&(���R���i�e����8�i���XW�P���Ɛ=����因��A�^c�3c8�E7�*l%ހ�1a���O���5FYL����}�/.LV��:�f�o=�>C���ͪ�����J�O��Hf�}E��w���[#/hoPPR61��䉍��^P�[ �Se59�n៤$
,C�u ��C���Є&V�p��x�ݔo�G������L�,nz]6F)�y�+=��в�iT�.@�3�%���
$�p�&O&U8�b�z���t���D��|�dA%(O_���0[�N���I�bs��@Ǵ�&���{ݫ��`���3�����4�":��h&�aAg��D�ڀ���k��� F�(#����+V�.o$ii�'���>	fS�SP��T}#�X�&�j�I7�@Z��i��*h�<�yB���ܵ��.jv��X��z�� <g��P�ҷ1��Rh﷬vI=�a���b�w�W�):^�<��u���$�P�,�sO�ϑ����0M�p�M���>��d�(����	��;�N"Bl�.i�Io�����<���a#qЈFjۉJ�v�a�&BC�p;�c��Ҽ�4�\Z	�Em�̯�>5b+/��NC�ݞ�[7�y��u�ڥk�j��o�g}�:��YIG6������@飯o�;NS�¤/,�'Gr��/ʵ]�CH�s.����!��t6�s#c��p8�S���$�E�Wz	\��D��w��׀�)nT"a��j���f;p�)Ga	���:w�,�?��M��t����C�투�ZB��b"�����@�F#��Y�s4:���r�>���9Dα�pFY�cNN߬X��Lx:��~��NP�E^�|c���HF��akk�qW�	(��HM?>9�ˑa�M���	B�tO����[w�I��Z��˶XA��`n�SaO����q�F�*9�xmo�^�ѳ=���8�ܪJ��JE�S��H;��:蓶 �
V����%���i�y���AF+)���۴��6��/"%��[¥6��F�~�3F��H!�y�q+�KF	�~��6zmpE�k����.��[�5�{���V*�:�R���f�T+Ob�ĉi�v �r��~�76r%C��9��a�ސ1d�v83VVAi.�COf��7��M�[��	���_��a�Of=L����k����ΏgYx*;�GX�I=E�M�E*��>;���u�ø�/��S@:�s,�-�e3,��yI�6q_	$�w�6r<�P�
1�����F�)�\�3��{	[�p��ÿ%�.�JZ�-���l>Y���zN/+�����������Op��ق���?L��kN�JӇ�T+.�@G����-C���=�{���M�j��%�l�cʗ*��`.�L?:%��X$d#0��� ��;�79�ׁNw�<2���J�%,��� o択+����H;��Xυ��-��|���w��'��C�������C+'��Ȅ�t�����c]t�6�[�p�2.a����SX�8�*�}G3�������<�e���	���S�{l m��{��7$:�+e	�t����t>���1�n��L.AĻ�2B���*c�)ߵd�P�7*2U@��J���t��G.*z�uAฝ��I*̲+���h�vt�b�0����g��$G�lAP���<8IZ��3w^v�ٞ��;͟��;�ޮ��$��S��d�9"�P�`��A2�����DEEE
�����!n,j���->/�f�+ʴ��叇�3�~�PpP�P�.d_�� �m�	j�{��e��ݨ��1ݪ��bܳ`9�>��O��jd�H�Ѩmp��K:����j�:-g�d��y�:�;�����ĞF�rv95�'UFF����&��
g1.j'6�D�j;�bT�eM~/j]����Yu[ܘ�āX��H��w;�!��|j���Y�.���2�[���\�����NT���oM�+>�#i�"�:�;6�:bI훭��wS����s>٥�c�#�|��2�
4��-oĠz�]����`9�g��i�>���D7}DT]��cR����_�l��s����N"GO�����68��;�"��۱�ͪ��S3J�[��$�Tn �EC�1ۢ.(@B���S�e\�E/�U���v�ɝh��Y��s�<��(2U�2}~��k��껇p�mƢ����1t�	��"#Q�؂�st���;*X��E5�S��_���{���23�6EGE�/��}8������:�.�D@va��T�f�o~@8i!&�h)9T��Rw4�[-�q��I�
�N�/O�y�A�"�F)��V�G S)��k���Zͤ�A� �q�yq'�%�˫mt�ِ����"5�
.G���Pb���
�2�<��^;������H*��y���*����l�i"��"O<a�� ��	cz�v�6�ބ㈲lbjt� s*}*�;5�&�2$8��&O/�j�)wTٯW�������"�s+�uK���d�;�2��A�����,)��/���m�]	��)�n�ΐ�v��9��ueC	i���'����_ʄv]�Y�����v�~��8�
K�
Dy���}�M]�=��rj$��-�|�jd���&�� �����.��t�@89(�IB���RJu"�逸�=mţ-/W��5�:E�.s<} �CN�B�-*b�����b,W�>��bق�C���y&pΑ��,�ٴ�}��Χ5��_��d�$��u����`Q0��,gۈIQ�XA�E��}���<�,ƹ���ѫt�F���^��|�Gx��8�Ȇ=^�l[A��U~Ēq%�YdD��_����3�ŗiƙW���vbp��Y��Kڮ�ji+tgy��*��q-�����	noo���ԟ�_��w��o��.�yj���ʉ2S8���Jj���֤a��e��E�d��
Y'z� �lt�g�fl�/���U�K�OVT��!�!�w���Jw6(G�r�;�tQ��������?��=�!cAf}�A�(�K]�xdf�Ņy� ��샇�#yn�W$2x�O�.6H�[�\ʪ)�JD{��b�順,5*ʃ3��y7��H��ġwsL�"y;pf��b�:s���lsc���f�c��[�W��n��XI�R�2.DՏ� �|�@�T������vz~D*�8KY��;�I*ː���E�$B
EY���W������'�㹓�v*}KY�;^�<�ZEW����b���;���c۬l%�-�؉��L��<�0�6X�go���Ԥ�e����rQ�)�C|��h_֜�Ls�m��@�f�F�X��j+��`�ɵ�<��uȏInb|��>���c����$A��S(μ���(���� �����t�~�<�u�*��B�T��I���~Tc��J7e�҉��Pe3�L���$��0��x�1
Bwم9<fx�E��S"m���Bvd=�a�}����� i0���*u97�'�c׏�,��)3��e��	� �eyl���F�p (�QK!�L{N�+Y?�l�֦l</kr0��g��lW��Pq1!�c��TB=Y�z�5��,ڞ4�n��=ԏ�ɛmp��~oJ���)�l|������>g�E��Ҙ�;�)�z��,,�cO������r_���O�g�B��m��l�f�'mi~�cŎx��.I
|cC���2P�`ǎ1�4�e��Ƣ��*�0&+yD���>��2�H�0MD��,��&�f,�rB �H�O��;t�9l�,w6���M%3��T��H��$�z��M��mC2���yY�4�*]Q��)���� ������G�wp�&�m�ȶ ������7����>K��D�C�&����˻����eI>n]��C��͖;v"����L.�J�*a@c���H>��A�8�������Js{��y��"��EY��ED����=6�c�R%�TC6�P��I�K��,N�.eJk���^��NW#j[a�!;e����5��iEj�D2�I�oO~��(�~R�5[���QJ��E��gR_ѷ�SݤP����:�^�~��>�Ez��CD�Z��:4��Apo2�H���J�-q�z��K)�{XQ�6ܶi�6�>������L�X"�]�/�x��1�G�#(�>R�r���<�0�S�&ͽ�p��χM^��r��t�Q�r�ͼ�l�jE׌G���l���Ǎ�-Dɨ�����w�#��6ʋ|QıcT�����v(���v��N��<�J�+P��_[^ۈX�u�u���]8݃�moo�4GU���T�j;��P#!���h�.�d�1u�J^�k���j�9ƠȮQ��D�VdBh3%�<�c�f>H��R��� Ȇurq]׀��<�i��*��M��w/���!>�©u�6���]\Uَ�L������X\��&�2���	[\���y�/�t�)"戇��3�>�a�T{,�;m�˰M�%�H�\�BC�]>"�1(�����a�o��nu<H��@����%��	�;�D-(�:�#] �a]nk�Y�[P���':��V�F!�I��%
T��Kt����*݌����I˘��4bn��K]���)�U��c�SͿ>����6���Fv�⬌���d���u�׼<�ѱ�$ō�i�1�M��@���=e¡����#���� ��q���i���{�W�E�^H82ސ�c�h�?>��)���[ ��fՖ���BU6��o�G�k�B���҆0����_d8�0���n��?���֐���w�V���)�������Au���C��&위�N-��?�\�n�T�^�4��ʕR	+ơ�A���e��V��m0�K`W�j��%
Oo ԅD��O
�&@��û�;(��������]\����9;s\>k+W������ĩ6;7'9̉ʦKFkN��2��BGƫ��:dY�j��J]u�������Ƴ��Ѷ�%�EX�y��)�����,:��n�&�O���B�� �}fprH���2ǩ+����B~�T9��[���pSʮ\���NX�����Z�������m�	�V��i�0�(wʈlk�;���:��~������]ި>�>d?���F�ءC�)'�C�ZMqn�o4Z�լW�c��E�e��nC�� ��Zn�3�Ec@>�+�dtjy�O������8D��Ƌ
)������:��m:í�S�0}>��!�/����O �J�hdo�~J����lM#��2�0T�"��X�P���,�¨�����9�����S��G�I.b`޲��	;svѮ^?g_|u���O_���/��m������Ǵ����q�.9��Q��@��~1�-���c笇���u~�7��B�I�m�O;��B�[/��2�"�+�/�I��a��)ٻk��
*����NY��
�gN�+�!��@�t�3��>\�@��=�s^�#Kg�weg�mf.��]��w{sͶ6�+���B�������˻�tn˳����K���pp҉E^�f
��q��C�/�Xf]�:�?<���Gn���=�j�J��I&�����h�.��S2���F����,D4i�.���wp��h����ve"�XmL�N�x;����&�WL�l�i���7�
�.�O
�k�l�
���!�g����hJR�c.!�vég<�����ꪞ�i���M����c3v��I�}��}��m�ӟo�7�޴;_\�+W.����6==�E�_[��Gx���B��,��!ԁ�z=��~g$>��������i�Q��򋝂<ZsbRC'D')�:��o��8��qn�cRd�GEw
s�s�`Am�5dWFxl�1��G�ؒ&'���?���M��ް��M����u��~9�����U*U�Y��;j��2P�?D�����:q�j�q���n�?�P��ƨ�?8�6m��)��P�m��eg!(D/��[�r�T)0>��Dj����=ɏ6=�@q��-���������6�Lp7��J}F����x�q��L�?Z�M�X��g2���I���Bh��Ľ��m��޷�'������7����K8����W�Ν�v��;q���΂�w����[E�\@���l��@����+�@(B����cR�(TM=�$�<��b�ԏa�y�?!����\��J�^���p�q���U$�*���? r��8�Pi<i ��C2	��s��;�?	��Ƹ?��vo~0C>��k��S��8m�s�C�k��mc��6lO�?/K�vzjʦ��A|ā?v�q����U��p�W��;�Ox�����Bu� נ��-�tf��<����2�QP��;7J�4�L��d��~]ǐH��	��]0~�KlR_�Ǥ�����ּ��#;��x=�q� ,CM��S�GQV�V�)�x��^6V�e|P3$�����Jt��K�Z�X�kDz�x+��%�Q�+|N�9�D�V�nd
Hk�],w֯)�R�o>>���SK��߈05�gXO�X���N���v��E�z��g����v�첝:u̎_��|�A��WW�Jݾ�^�2rx#J����hƯK�,Ê�.��a�b�k�͹����!�+�-q(G#�Y�*ļ�������.˔=�곒W���-6�OHC��c��h߉J{j-[��]� v��?DY�FUo�f�~��)����'���N��%�7����2�k�+mP��*#�S��Ib�h�#��� �����uY��+7�����j�
]��M(�����F��f�'��ۅ�gt3�"�3�����)��|w�z?9ƅ�����Cn%�!!��yy��1N��T{f�׳��2f�0��e�._�,��fnFv�W;�U�?��6A��fA��<Z�� 4؆کl鍌C�w�u�N�y��F��6(��6�<�����q̍\�Ęe5I��2q�M٨'����<�x�/��s$�3�|Z^i�B��*��1r�^�:?dj�ι�$Ɲ�M�r�H�W�Q�9���A�����;��C"\^�I�u��6�JF6RG�[���E��W�7Dq��w���}�]J�ҊRDK��^����br��5��_'����$'p5��Eo������p\o�X����e_�n\�l�N,��̔����n���<��-u\o�d<����Č���U��i��2��c����]4�7�176)E
9V�vp^G��T�Y�G������r�J�����)Q�s�,QIF}�hG50�VS��6�h��#Bz�h�?|t&��q폅��n.�O�5y�B5�U�u!�i"�IJ�������R��D����m9u��Nc�iبqR��%�̔�L??�����M}�C��T��ܦ�G"����m{���ͼD�#I��zc��z�5���BE.��g��	�#�m���cKs��rξ�����?m�~s�nߺf�.����`�a�Y}�c)��`�ڢ�,o�#�Q�|Ջ�Q��9,[s�Cf��b���<䷉�����=�Ww|~�y��6u'��~�|��צ���t
�����z���.}\7���ۢh�FA��zR�z�hg�4�vb,�l#���g�%��T��pps%�EL�/�$���Q�a�[��nRp�����Q��i���U8���+�}ԭ���Qu�g�<���ğq��qmj�1t�#x��[��X�8��-'��'CGJ�v!�9��|�cE��\��'�(ml$d��Q�)��äD�Q�+gWF�ŕ��?_����y��m˱={zٮ_�d�|uǾ���ݼ~�.�;c��m
�N�Xث��A�l}mC'2h���Cu��>�xbT���@=�q��B}�$��q�������"�+""����ľ�C_�r�W�r�,��1#ʦ]��UQ�5��; �C������N}����~0(_�Q�	8&�$wf\�ۮ!UBV��Bi���]�_Ҋz�%?ORN�i��[m�R~�X��K�V߸Sړ
[T���YqE��(�#�i	��+�}�Α7���	!m*]]?�R�G����vo�I��3gNصk�/�؟��n���}��M���u��r���p��#��]P㄰��_6�ۀZ�莒�y�@Q�_H�Q^Ar"-�F����R .�U�R[6M6�:7�j�p^�Q�"(_�T@�����z��T�`�R[�y�u��+�*���P�����7�̉vB(;�\�F6�e�eh�y*���\lOg|
�m\���p"�Ɇ>���fEYl�G:
A��KΨ�n���� 0@Ͽ�i�D��k�?*ܦ솺��@��#���G&p��vw�/Q^���&ٮ��o\_�����O��g,�_���v|i�fg�������>�����#�{��mmnʖ���i�Rn�B���bh�.2��L@�uz���w�8V<T�t!��S�m>���'~w��6�w����cRYO��s�u N����⬭\>o�o]�;����_\���U��w��O��7_ݶsgOb��Z�m�X�yWNN�	::&��Udy�W	�˨�Z�9���g/��
r娺ӊPw�W�%%���"���C��Á����9�����~�Ywٹ1_[�*���b9��'���tl`z��I��3K�""�}�ǂ�j:ȁ��A�#"�U�r���9yxr!e:�:�����=�tJ������v��i�y�
��v�ʊ]8w֎�c;�c�펽|�f���c���d�޼��6���Ol���'���yG���ۯD
�>���� ���>�w��~3
M*?&��9i��&r�G�#�9�8�L�'zp����k��U�N��\�����>�h�N/���'�ڕ�v��e��Wl��y;u������Lz��ԉ-�8~�����r�1���+�n�M�b�,��ЦcJ}���_�*���O��?:4�q�	�8͋�|�=��!BQ�Lw	kƮ�i�czn��nI���;��P��܈7��4��9�� -Է$t=������ӂ��vtD�8Ru��-@{m�@� y�ȕ���h6�������X��ɱ�u�]Y�hǖ��	�L�[[����&ڧ��O��׻�ړG�m��{=�@�M���|�4{�>ϯÂu�6
[�;,O����=�]����y��S0�X������ޝ6u��kM�xTwlD8Q�9���s�̅�FD��K:f�<�x�ѷo�a�c<T6l�������A���v��q�~��ݼ~ٮ^�dgϜ���E�:�(���q�8˚�L�@)�(P{�Q?;EX����@��,��đ[W[��d�4]���AE��u�Y���3�g��sNJp84$��|����;�
�������ۅ��0F�� '���8u�9��~V@��C����>1��2�Z��P^�.�QP��^jJtӨT:Q#�&�]������ٳ���؞��7/˹�t���������c���+����7��Ϗ��݇���k[[]Ǣ�?r�/����$�Z�:��?�.�d��o]�
��f���12����]�{Eݵ�g�z�S�HqEK^�j���zIz�;G�x��3�¡uJY���*�i�'��dkp�
��30ċ�j yDꤦ�Ot~"<z��v ����Q:��@��v�u��!�7V1�,�3���i�����w�mcck�ߐ�����Y�pn�nݸd_ܹf�n^������4d������Q/m�/�T������B�ԇ�^����,��F�=���Ϲu ��뎭���	;4���
t�q^ԥ0:�^:
l��RM��Q�ׄ��Ԥ��7]�ea��HM�h:Z�A�9A%�U�P_Q
J�R���q�P�t �Y+� �2�������I:28Q �D��߱UMcU�j*�s�z]����1��ʯ�;6c׮�����n_�oE8�|L�f�׼�����m���c�������믏m}}�98���4ɇ�A����l[w�]��v�[c���!�i���j"R��W:w���� �~K���@���Ȯv�EZ�\�
�bצ؈A�'f yFP�[�ƕ%�<ϭ%?Ì��;挷���FUW6h@Nq��0dS�Qr���!�C��!��|,a,X/����x$Q&�g�?����kֆ�����2�(���Nʑ�\߰g�_��'/���5[�������=�����^���-�����ܹjǖ�����2�����Ϭƺ�|*�r�#�W�%���P�aX��Ƶ&�[:�(w;gIGU�b*Qa���V�S�O�n��kZy�tsu�V:��E.���
4�1�|/k�J7�������㤝�]���E�t!.����p`�3(��$��@.@�rZ��*yn�B���ϯB����&�ю�^vPq���g|B��C~��F=-��r\'�:�TMT�e�, :5_CxYw?��JuW�	Y�Q�y��P}ht�neB�=���Q�vj�*��Q�ZNF�u�� ذ~W�1���vsr�=�[rl�f��c�v��	�⋫���kv��e;��-����$����b9����xz`?�}d/_�bzс���D�O�پΗ���-I��3�nT�4e��{��d�<�Z�.W/,S!�~��֕�^/�*Jq�h����ady��(®��,���V��^��f%��a��q6F�e	�"��%!��-���h���@E�pI��|D�m�P-�r�!� r�dHd!?j���t����'!ɗ���a�&�+5���G�\��&Y ��\?�\�ʼ8�|�y�ڊ��=�f���R�]�td�����HET\ʊ���\�z*o�3ɨ�{X��P�
2XO~?�ı�X��5�m�W�q�a��\�w������9[XX������4	Ux3lvf�f��l~~N�76���6�;�G�x�����v7�K!ļ\']+ �Y��)i���E
^�L<^�� ���׌j���W�C@}���A�
\���Z̵a�	 ��\X�*c����s{�J P>}�ӑV$�CU/{�S�������C�G9<W�#�]Dt9⍍L.+��z���q�t90ɝ�1�v��9����}��I[Z�s�K6u����յm��[�dN疕+��I�V���b��O� :)al*\&u�� ��RY�An�Ri�G��u�`�U��R����39	��AB��h�-Á�Q���.�Y�L����,mC����_�ɴ��@�'���vQ�rn�O~��:N(M�zJ4�J_��V�\�(cg�ŉ6`=�'R��x����|��*�`�e�Ǧ���2�����oo��W�̩�pl��-�2ܷ���/��׿>��������C8�X9Vh?�[4,=��3\h_�"�I� ������K&8��V� %�����EVal�uP��?�C:/(A���l긞jFĸS"�xʱW�kQ���a'1C��"��X�޲m1��CFE>��
c�6H�/���:U>ǽ�y�+�.d�~�Sn}e$/���&��A� ��!{��?�u��$y�*�h��S�S�xZcd�� "N�ΊP�9�3(��Ԗ\��l���I�����P��A}��V��Ey��� ��f�P�X�e�T�sC&eG9�u��y���/��>d՚�8W�rcȲ"�����~�me_�����h\�SE\���*D<���N�/�� L�i��S��7O��m��87��-��,�f�m/��3�Ņi8��r~i���5к����ܬ��>�˛Gt|i;�cL��i�o�-u*!l�E�,W����B�vnf�Ћg�,D4޴Ə7�4OT�|1?x�)T�
(B��$�{��:����
YI���.zH�'Q��<�L�/ӱ%%�,��:	��<�*d]�#D�9�rN���B�Z����O�������/�ԗ@�8�]����]��	��2�Y:��s�έI�R�LK9Pvq?Q�o$��e����8>�(�wG������8޹��S��,=ރHGSm�~ܹ���U�����Υs��������(�<ʕ���6z{Nl#��%��$lQvI%�B')(�*R3TiE��n`}��/XV�)��5-���~�����xWK�v��1�}���+z�oEX�_�i8�{����go�n�Ç��o߿ =��s��pҎ3��pn���ґ��0�ぐ�F�X��H������tec.�����=
�ض�[��4�	��	�|1 ���y���	C�:�үV�yN[R�69�-�-j!�P0�񪞷�
��l�W��'&ٍ]�����Ӏ��R~ ��q]Q�s�.j�آ�G�-�e Kj���렝d�b*��5��(�`8�ì��N�� ���CB�~<�Ě<E/�7�sk!x�[���T֭z�L�4�Pʕ̰ɐ\o�˝G�/�#��Fv/W��#��]Bu(��YT���Ნɣ�]�V�|��*]�8��䴯�ZG�����|���#��NOÉ��;����1���<��eӛ����e���'�Y�ɱ��Z��+���PYU^ 盃�&�Z^��_TO9�<�eyٔ�W��B:+��(�}HuX7�3DTs���.����ַ�]���/Ҿ�O?��k[�z<Ւ?dQ9� �J#IY"?�
u�`o�uMy���ώЛ���C���. =��t>��2$8ut#�Vwn�4u����?����N��tEԼ�
����W)N���ΰWL�QPe �#SR��y��˯0�  ����-(,͹��y��g���W:�����A(����yY/��@|�Nb��)�2���ύq���&L�u��H'?T��5�:���\�6o�F��%��4�B�J���z��*{z�����@��_Uam����:�����잝;s̮_;o�|uC���[8�3�S{�X��^�ڶ�?��������_��/�>�ׯW�p�=��H�*�=�kd�U������thsG4�X��q�)³nZ	�mùM�>O����t��Q!�<�����U��I� �}��PǪ�b���G^T��u�G��W��o !��U�����2N�Y(�ҙ�tL���鱔[ɣ�\�)�1�Tֆ�S�.td[=�l�"�yl��]����<]G���2֕��]`��7�AU��$d�����j)�B&#l��5�FGD�Bg�B�C3�L�2*� �Y���i���ϼѣs>��g=��8U�\��wq)�6���]]��/*m�|��=У
;|�x���[t�r�f���=$�����M
��^�Q��@�%_٘Ϗ���`�j���®\�1P��`Q��X�E\��`=�?خqn#/�ƈi��!�*	㨁�6R��ENS�`Vɑ���tbS9d�0$R�<޲6�D.�9W`�J'������O�cZ�&��+��i��tn�X���%��Y����rRՄm���k��x+�%B�E�D�4;Ec�ÜU,J]�G�R�e^��R�}�_�1O�l���g���hteTi���x�@�c��*���5U��Ɛ_Oq��3���OO�aq��v��{Ӧ_Z����O������%;w��-�cr������}��}=|c�����o��>���`��`.ltnyկF�\�1�0h�2���+�"=��,�DG@� �M��K�ƹ�Y���#67���vCyI�>|��>]�����������ֈ��
�
�|��ykfk�t����6~k4yF��h��A
��P��3<�紆���O��3�F[ĝj��6��A�
�E8��p
��I��͇�����5�d�����_���'o���m�-
�5;7e'O.إ���\~���r�N��ci�e���#�1��}�')�;��f@�-�w�R�q8��m�i�K�u��
��H���#w��,�ôU��\Β�;���۩>�;�^+�B���P�*� M�j����'�&��L���9YA|��������e�D�>�G����lR�\�b=���,��;�Rd5W;��AW<�Dq7�.��tĳ{N\\"?�D��C� ��W�r<,�G��l�Ε5�Lz�8��U�����*{pj;\���O���`��������Ν�/����]�r�I8�s�8e�p��o���{��㱿��,���������cӳ� �K��E L�Յ�,Pʈ�yI7Ȭ��3&�+����ؕP�sk�MA��~�`5g	~��Q!��1�oc�?c�u2�È��N�&�X���>��_��Q���?
%���Q�O�;i3������F%�{]�j�64��tP6d��'���^x�x>�OY�VY���y��z~�-����"�,V��*����
\:���'�92Q�Q?���`��.5���L��G�<x��d	��N|N��P5�����t�_�����mml��ښmm��;nhhnv�fg���#���;�y�laq^��mv��o����m"�x�.��:�l�u��7�8�C�Q���u�C"�*������h�Y�"na�(%�]�v9?1��z�V��+��6X�wm��lO]�Y%��4�I�����;�ȐN�Y3j�.r�c0L}����YU���/���1uCG��<�l��"�i�ܧ�ݹ=ѽsϾ���)d<C�8Pim�J�"o(?�V����Mn�\Q�;N�\���VmE=e���cȴ�7u�����rT��\$��F�cQDb'Rn�x_�C�.�R*�3���*������;�;�{[�;X�<Y�´mǎM�*��]��bׯ_�U�%;����n̴۷�w�ѓ���OO�ؽ�O�ŋ7X�pQ{��"�F-������MEP\4xq�9�H�SЕ��<PE��ӥ��C9ntq�CQ�j�"��A�����Q�S�]��s�h���п��tM����rj�:��'JP ���G��u�H��]�C�͂�/y���T (29��+�B䋘�ۧ�kި �G+��.����t@�ݛ�S;�7�W����������{���ӷ���������ٹ;}�]�|�n�Ĺ��%;w�[��ys4~�B5��@��,��R5_���媫+��(w���q2��G��O�f�#Vϝ��/���ޯn����p&� 8�
��:h�V��QN>8)y�ԝ$R\	�Yp�9*ā�g\wt� <|�S��O9,��PW���!#��_BP3��&�{��i?x@�(�z�-l~B��I�MfgUrXڀy�P�ʛ��W��=,y$7�$��L�����MtӰ���x\���G�q����_0b�`}����ރwۖ�������7���؝;7��y>�0��Ե�,��pl����?�O?=��/���3|wnN>$�6�?۰},��*T�Pq��"/}�d)��H�q�uM����&� B�g�WJ8_c~�Nb�PPq�#-�����:0n��t2TwDufK~�0�*&��a�|BfS�ِ�~`�9��O�+h��,��a}���|R)UsOcT�����^��*�cg�$xG�H�)谶�:�~LeoX_uH�GcQސg�Xq�q�O�i+��P���-dQ���|ʊh���A�����Ԋ[�y���x���N�/�>��=LF�E��(@t�΀��s�u�F���
��3q�
�旮X�gfp����-�����@o^�qyg�o��I�w�w��B�ٸ�}��Y�S��=�}Ɣ́��`Ȳ�>x��-�a1tEb_1�r������Jn��6?(�w*�e���v��1>����.ʨ,�Dv����9l$�RpJc"�@�<g�r��$(�p2�H���:�<B����	뢶Tpø�톢�j)v�IF��d���&&�'&��P�pn���a}VQ]V&�"��M�3�ި��C���`9J�-Vu�H#��N�=��qd<5>���6?���	8��{��4?eΟ���W��n����]�xΎ[��m�
����?yo?������G����ɓ�X��Y8����#��}��gΉ2�S?�3�G���2��S�Nur�*�7��*�*JOD㑙�2�ҝ�l(
��%�ǚ~���<ױ�v�c�-gEQ����9/�b�:���z8M�W3P���U�!�,�x|�h�g�T!?J{���r{���HDRصG�k6�lW�u�!98��+������g�*U�+m��h% ��C��b�&R���E��|�S2��&�i�G�İ�C�m�����y�A9���sd��B�QL���2��UQ0��BiK���_�!�����ɾGt�wZ��� �Ga�3�Y���4��s�(��w��p���#�8��WD�;p�y�ͱ�F)�QEǢe��P��o���X-�I��ͩE���pQj�ho�����&���/�N$�����ӥ=fɯ��E��v�ȧ��ܒ��0bN0Yέ�c}���-"^Er\'vFz����^���un�r)�yrn�PF=��۵-���32�Q9��@����/O⮐�m��[&��(�Q�(���c��W������2XAvN��q  �4���c�`M^� .ó>�~).�ԉ�� �G~eC~|d\� �S�j	�D^�]���"��f$J�7uGn�����t�����8&\dh�)L��pjr�Bڱi��g'���v��5��˛�����k]>��ŌN��m���w��ߟ�_�rOwl�=}���8��6=�)8�Ё���nm��ւ�St�O&�!��0�����Qԡx�q:@P����r���m�Kcy2J4t-��'2^*9�4��Sv����H���~�BX���R�F+Mt�9aW�"�5��AP�m���6,� �=���@��:��Ou�W���j�FN��� �y-�	EJ麜�t@c�9��Q���!̈́들�ev�VF3���rɯx%���s$�D��y�s��3�y�����O��Lօ�����/F(��g��j��"o�a;���|j�aCD�1pA�S�O*�|l<'��O�9���.��+I��oǏ-¹�����߲��W�k����C�xc}���O{���M-:I�	�uu'�����Y�s���7ϭ�"��]#��Ԛ3#Q�$���&dIP����6u� 'R�t�h?�$"�#9��<�lzũ�[�[�O�B�� "A��t�GB�ewl%K�i�A��L�(]C_�S�,l��r��7�S!ۛ��g�;tn�0�&��[:�� ��(Ty�&ƎkB1��d)��"�3�!�c!�. E�V~ʓL�]��/� +�)�gǘ��1�����P<�*���TQ��w�6��V��OU�ktӽ K�	�}�B��x)ʈa7l�9g->���m9�z���6�?�c;i��,۵+��ͫz�������E��j���kumמ>]�~xj��}=g����u��/�^l�N0�Mٲ-�>��0mYu���Ucΐi�z�L�� ]�r���$��ʦ9\�W�F@Dҩ+��ȹ�����#�S�:�]X�]Uu�m��^�Y�)�{�n�}�,�TC���'�:�~v;SlU�s �,tBhҽ�2�B����6�y��D�?��a�9/9��&�K>��ѐ
��܃RTdf�Y/<��F/2�&f�����,���9c�d�%UŇ�;,���{��w)j���z�o<��\ޤ�ٛ�w�7�ٳ����'�'��؛������wo'l�ج]^9i�n\�[7/���8��3�k�ۛ��������?��@�j�5
�VW���Q�r�y-��f���XT�!G{ű1�mx�|1UP�;��H�*YV
�4ɩ
UKyQ�� [�q�Ǟ2��+�����$���VT�U��$�H**i�m���f{��z�����\8M�
�M#�n2=�r���<66�8�tR���		�h?�~(�}���,I�k�����h�H����N�qӤ`�ONf�NAd������m�H\����d_~q�n����0?Fw%ױ�=y�e?��FoE��ow�уg���:�q����c�y����&!@�;D�M��tH�r�Bo(�q��C6u�)Յ�� Ac��x��9I.��@Hg=6��U�O��?�1�Q��;'b��+uh��f��윥]"����>��r2~�U���\���>���X�2�"X0�A�9?�<�.�]��D��1�]�#Ue�2R�.��2��!�
R�bfz\wj�5eŴqMc
"պ�,�ѐƐ. ��(ў�����*�i���மoړ'/��{O���^��z6��bI����������e9�7�]�s�����m��9�ZL��M9(���W���< �#�(#��X!�_���?E�G��Դ�=U�*��|]��m�9��� Fr ����T;< �'1��4)])�]��X��Sn��}pr�4`MyU�q6�0����k�2�s;O���N��|�JՈ(�M�S�lۓ:y��p	ا�"D���� F�-aw�bbK�sv��I�~u���t���\>�;��������V��÷v���v��3{�������|��3657�NB6[��C[�1��N�����;�N夌x���V�܆r5?��{��P����u�H���v�?N��C��:Q0c9��ƿ��+�#�0����(�n(�&^Ѷ҉�yk>T(�u�P���&|,j���8�Aٵ �T9�N)ꓣ�H�M򴏋8�XA����� Ƅ�����^�p��os�#tޝ��߾߰'O_��_�� ��޾ݴ>�ƿ�=sr�._:i׮������y�Aaa֦���Q��A��b�T�;6�c�o#�T�M'2Ty�� ����C��;E~[�CT�	�ǯ�=ߏ�(^��ϊh����U֋X?��*U�З�ܒ�[�"�o8����щb@�BgF�uD��Q0�2�/唆	
�"��:^Q�W7p7�|Z���N-�Vɰ^S�Y���:mv�p�a��w}����p�xw{�ڞ-��ڹ3���;��/���K�6���༮����Z�~���޼Z����M�����hަ�u��&��Mұ�U4rI�!+h���6�x'J�J�+�VL�_ē@\��ٽiÉ?Ћ��°��K��.�����Ѧ��",��e�B�6��=�<ҾҲ2w��}폣u^�L�N�{��&�-���v-6�[K@�W�	�u9~:I�\��E��o �Y��U��P_�r=�5a�>T���v�T���(��3�N-É}���7��TP�`�sM��o�a|��c'�����;m|�����rl������3{��ml�U�`�r�Sv��"ۓ���Kv��E�p�-���\�e�k�yC��7m�[�O6H��xJ������<���u3�K!f��&����q�HFH��&Z�f�55\?�p]�z��a����b^#p4��X�JY�qTX1J�J}y��B^,�BL������4ª��D�r�3$�q'm��v2?�N���NC����Ⱦ����V9�4Td���OT|3'2�{L:�3v��]Y�hׯ��ʅsv�Բ��.,*������={o�_y����!��5gy�"�87Й�3�������.�x��1F>��Ԯ������<��B=����8��u5���!U�j͝O�ZmΖ9�2�P�Ie�
箎_UgYM� �����@c���$��D����O���c2��q�zE^�r����ڄ��zP3i''�
�@4����.CRe�E��!O�ﱅ�+'W�<���Lht�X(�2?o��Ĵބ���[=����>�/�l}c`�pX�c�cK3v��1=��ŝ�v����g`;[�{�9���	��a�ãB����o��Ic�BW���r�]Q�{���3��w��2�lsD���E=έ�{g�T�`D�RK��و�"�Ӟ��?���kAP�F�@��L���St>S��ʓC�+��.���?��H`�_��T�Ԕ��@s��@Ԥ�O�Aa�b��$�VN-B�7���GT��U��w� ܱ��	8�����v��uݵ=s�-�J����q�X߼ݴ��>���v�����^�x��	8��">��?������ǘ��}��r,�64v�
�:��j
e\��I%e��&�Nd~�lF�6
{A��R��kUL�:��ء���E��(	s���?��y
q7��tqJ�����0�B����:=У`�j�0I�^:��)��QU+��_�M*p��� ��Ʈo����+�î込>��R�u��p�B�k�*����L;�6
n���]h�ЦS��V�)��!�T˧�RޑB`��*��7��,ob��:kk�z3_�������}�o��3.�|��y�~�}��8�����)����y`��������+�Đ�1?�{��nS�)@�P1U=*:z�Q@��L�x��ۓ%�q��Ne����>W7�)X�AW��;?J���çE-����+2.x�ź ��\5w`�d5��(�#�Q�D�NJM^�uo
h�Pm�-j:K�#u������O%A
�q񕬐�f�d����K���s�DX(��L��J��"Z#��v�A��prp��˳��Qo�#D�t��2=�I��l�,��\^Կ��_7n���Kg�ر8��8QN�����<ygw�>�c{�����^�|g�\ȰX�o|��|���`�m����bT�\#����B�ϸ�����	%'�+�Îe,5w<�uS`NA�a�y��4���w�E�(4�R�UE�4�ꦗ�b$��N��",2�!���Ơ�&����ǽ�� �e!=�Pu�Z�W�ҥ�Q��j�aDSu=�Q:=��96	���Oö�ݦ~}��3_��vʨ��i��4��{��z�V�*�>����%_#�3�+�ty�s��a������Z�5���	�tN=j0/ڊsJ�l�z",P^�Jf���\�����)�-T����]/f�]��΄���}��<xf��?�'��������c�la~�N�Z�8��o_�[�."~�N��_��ƻ�?�I1�8��-:���]�g>,��r�@��o�U��sb�EO����c0�#�q�:�Q�ėH���"m��2�W������gG!�R��\�;���������U������H�5�*;�d���䙺�տ~���8=� g�&���|<D�X8��zS����tx��r!.�CI.���� ����;P������2��#���(�����z;8 p�I9W(RU��x"uB�3e��
X}��Щ&ڀ/����ضl�D�x�A�cKQ~E9�"P�(�0M��oB_����9���b���x�J�;���q����ϭ�U�����]�z���������v��Y-H3�S0��~@������_��o��_��W{�蕞����S�)F�\�4P�y�ƄN���Ƙ�D��,ט�(!�+(ŒO/#g�X���:�9�n�A��BD´qn�H�'���P������!���c�O7�a�E��NCR���>A��kd{ߝ����.���m�<ȁ,�~"� ���La! |��u�uN�z� ��Ff��y�5z�l� )1Ƶ�:-V�G%�\�_��0@��N�j���u@�X��gV�V�Ћ��|�B\R�D}Pqm�����7\bt�7`�
41ƽ��6���Mا�U	䱍���+�<E�����D6�9�����,�z���`�F,�N�/%���5D�(�|�����X�P����5�2��l��|�,�����1�$��B��\�����#���8�0��"�F(�u��}�)��.�6h�)����aڎ-��x�-�����tNѷ�ض���g��S����1�Ќ�&�O��C��?tw}��B�z����'�J���M���ڻ��x�9�5�L~׼C(��UD�뉘�)�9����h�p�B&e�Z���eVB8�CN>�̀�2�sJe����)�B���ؠ��$9�r2_�a|��\�����������k_��wk��[�s��(�(GP*�B��!��CF��y�K9�/R�$����9� ��}t���m=�x�y�@�:�>pn���p��t�*��t�,��/�����b�FIe�c�l�<<�Vu��*e�|P�z�?/ggu�O5ן`0�i���~%����#&��Ζm���٩=�xWշ�؟����ڞ<�`s���s��x���"���q����C{�+���71v�z�;�l�[���it"�xc�b�A;E4�/��n_��2������[�:.��d)Oj�	��L>ƪ[Q�{��M��A6�a����'��X��C'�ŁUkP;�t��
2o2A��<n2T�*tDP:��KD2XDB�Phx�&<_�-�~j^�����L)+�DY72LD{C��l�*��wu��jy�ۤ/��5<����a��|��M4�D��E�3"�j��1+��V��*����ꗚ��r�a@�ܪ�Y7�)~��z����C�J��[�^'�|������p���2^@�드p䢂�Kq�)��G����|�K^p�vʵڋ�K���cJY�3�&U��a;��h�G�,��|�p����t<==ess�G���;|�(��s��� ��6N�t\��~�=�#�������t �2�T�0R�m(�F��/���?e��a�n��YI�njīR��^��x,K�ґ�E�i�ךg��RF#=��b�0wl�E�`�/�ʔ�g�a��s�6�3�h�?�vlq�ΜZ������ml���]p�DYA��s�T��Ƃ�ܩ�snU�
R����4
9��:]��ҧ��`��il��/P���@}�� ��8I��Jy����Duډ�e���RBB�j�"����(��i�:�\c�r��&(��i]�C�	8��OL�y�-l��`�-/���W��;��֭�v��q]]���ξ�x�f�������{8����c��������x���R�MG���n��Qݻ�]��ު�$�sW�"�{���r���Ni�k��ݠ3͈��%B��;:�.��M��`e�{�.ɂL����g �6�5���F��=u��a�=�Oĝ7B)#.V�Y�B=��i�1�u1��N�Cԉ��
�8��ه�P;�@� ���Z�:>uC������1&��s�]~��m/g?x6�K��4e�<QL�
�RR�9<ҩ��d� �@�S_�|�`W�.�x�\�� ,"rf[s�� �e�k�
��x�T���S5�3r,���ֳ�{X��լ�������GY�����b�.��H~� l���KwW����a[�M�����́���x�ҹ]X\���E�jV���;[]}�s
�
���N0l����$��3�a��	ŋ��A��5��A�m�x�V�'Z�H����Ƥ�����mv�MH̒/��I�F�^.y�J'���r��#d=�J:��)E�X�c�:�.Ǥ�� ���4��I��Um���Q�}����B)�Q�����d�^ ����Y�f����:R��C�U|��u��q�>}��ѕ�e5���Mms�����@-4޿8�jt�r�!�έcBN��������;�����!�x��Ec����pt�~؉v��)�q��d�h'O.��;��Q��7����k��G�#ܧO���58�8nx�]�`��h�,v�ŏ�]Q�����>���l�����$���[?ب��E�=up�M@z��[\�;�b]!�9V���_��Ar�B���ᐵ>)g�<v���wز�?H���y��U����Ď�&�J��E=����N�9��GD��o��`�ˎ��Q���g��r�ynڏ�� ˺�Ҿ���e�͜*��e7��_��yY��1'a��qL$B�~�W�V����8��-��|ݴ`=��N�~����e��ti	b<����X_�<emO����~&[�Ue'��7�����-{�s�O?=�9�=x��^�Z��-���6[\��N��s޾��
��<�2����-���5���ُ�S�b�}����[>d�.��+F�|��Դy~ۦЋ��B�����f�~<9}���К�p�8��lRP7iv����#�o ��lɟ�<R���(G�6Tv�&_T���$FT~F����Z>��E��}�*u����vn�N�Z�[�V��oo�nܼl���p�j���m������9�����X�8�f�<��,|K:���v��bD�z����}�wu��]Q;(*BAa0Hà!��A�ps�AgmC�vz���N��A�pr��u�*�f�qŚ��V�ٔ�-)�E�/'X�K��<*�P��2G6Y�:�{�F[PW��~�Q��|��(��>[a״��"���;��5}2��
r*�)5
ԡ��t�mu��$����&��p*o�܈�肼�̑�Р��SY�!��C�W��"�g����|��&.��!��!W�4��d]����|.����rx��䷜֤thIX�����ɥ�Z�*Sy��>|x�ڻ�;e�k;����w�9�����[�;o�P��	����S���ƍ�v���x�[�����m���`k`{;�ON.H� K@����rp�j�9sG�o�=یy����lrh1��;��Z��Qf�ڋ�
�_Ą`#�z�I}v�*ZC*�^��a,$�x�;�\t�:8�b��1�����ע> ���&}~Ѹ��[ �9���є�Ưܹ�nc�ل�[H���y�.�?i_}u���v���9���٢3\���X���>���>�G��؛7�w���ﲝ���s�n����ҙ�~��eI�f�L�a���$|0I���DwJϓ/ Ht����-����5��P<l���i�mNN>`�`��*R窰���(��� ��e����fX��P���%�j��DC?�V��XSY�K|k"S���-M�X}��x#��\�D�O#rc�Ea�,ۖ�<,\dC��oه~"K��"ԗ�����Z�����\���Z�it!�$,��)+w\Q��q9�q'B� 7]'_�Q��Z�w�X�s���(��l��X�'flwg�VW���=|��=~m/_����\�T�7df��3Kv��	[Y9mgq���(�c2���x�&M���oRc�?0�c�����Aj��@:�J��S�6LiQ�a$/���1U�3 #�:�)��;�;A�LT��x�[�Yd�x#��.�8p����A��>$d	]6�Dc��8�2�t�󽁶�ɷc~Gyp�v����cr����sv��y��?e���=}������mn���W����+��Gv�ק��=�V��zƦ�G�yMb�����kN{�����#�I����іi�s�Ȉg���y<���Ƃ�(.r�d�����6l����{�� ���~5�;޾���;�����BPn�T���SuȲ%��CD�5��F 4muJ��]��oR5�PT�c,q�+�r�Ť�mM�F�W����G�L��w���Ev%�S��h�Dؕ�i�M-��U9��h��6�z$�a��O��狒�;|��u:H�9W5�����|��Swfݩ�����rwU�s�e�?p2���i����kH| ��j�e[��^9oU�P%��r�!Estn���mjf*�����Q���=z�V�-�[$;��;�<gW���˗�㼴�gs�n7�_���Z`�]�w����zt���>3�X�F�1�:���/Ͽj�?0��}0Eal�qQ���J�A�W'�S��S�"���D;���O��@�j!��v�o���4���.3}rDP�*I��-��ǃ�ٌә�ן�|�{8�]�/���1���_�ˁ�:I�`�سc����)�v��]�v�.^<c�K��b\�7�vp��f����Ǐ_ً��mk���r[�d��=��h橃8���6�j6%©ʗ;}:�сŒ�at�z�݋}�c�S��i'�5��3@�~��	H!l*�؉hs�+1�F!;4�Us�<_Dc����VMZ��rsv�(w@r[�T��q�R��)�Ac^�u�E:"٢�}J�!����(��1��x�Ǖ��}��e�� �EH���"Q���+�n���].���6�����|XdG�?�
*��m� �0�Z�O�]��%	JB%���8�K'J��a:�tl�v�mg���`=��E�$��k7d�G=��oR�S�6���x>8A~U��$P7����2�?ǹdjζ8w��pn��e|u��w�pp�lr��4N)������9�q��� �?b��FM\ �ݷtx��e��G����������u�Q�
AZ�h+���G�:5�dnHI�pW�zT��*��Î�&�i���2'�?A�Gݬ�ǑB�oJ]��&f�We���`R2{)�L,��1u���;�=ߋ�w˪ࢨ���.N��d����ڔ?؎��8C�+�Q����`��������P�(�eI/���,�^��#��4�J$��>�Ni�~�.Q�����j��ͅ)d;���hΈ2�e��Pl�<(��2��ٔ��r�-�=��-�Pje�e;;X ���٥Kg�8����Uė�-`.������l�/�_ٯ�>�{�_�۷���w"� �m�rq�b̯�y�R��\�j�FQvW��c��%a�v~ȗ�Rq@6G�g�c�;�rl��1���Q�=xB�C��1mv��읖,�8�>�"��r�P?�t�D�9�c�)�=jx��:�_y<���;�] �:4����t ��j��>�-�I^�M��L]A)�I��܀kD� ��d�B�(̴����3�-�R���H�RE#�g�6�:���B�7��T�("u��r����%����<y\���~���A��6��`���Q�Wp�.�+c���uI|����yNuH}+��%BիC�=^.'��-�!>_������_��v�&tr��w�d�օ�̧xnh �,m7D��x����l�?B	�4��P�H�&30�*�X�znm�	X_�/~�x|y���lq:�ש��Y�[���ݳ�` �x�sۚ����2r}ْ�a�!���K�`v���PD�Z��<?��#8���Y�:~�(�Z���!��ȧ!!�eA��� �µ��+ç�8�D9�P�\Ĵ(�"Qe�N�JG"�`�8��I������Ev��{����Vk�e�u��W5,՘���߼�y����Au[\���'��d*�{n��K��"��JCT����C�g��]�T}�P�s��%�%B�(��4끢�����<�`�W)%!?�ȫ)�M� $bx9���[���7:w�xG`sp���'�ԩ%�x�]�zN�Y[\��(���E��Wk���{���uf}���݁W�X��\���O�P���TRV�H\
����B-�\ȩ#��©5�{m�;Xhw���'��ܹe[Y9cW����g�$�4\uA��h�c^8�_������(�D.�N"*F]���[���}N�c���������fK�� ����6j��)2�<�{3f<�/�v��A�Q�R{Q�i�uD�[���@]�%��8����M��g_�ä=vC㠆�ʊh+�p%"D��;r�����g����=L�g���h����*=`S:���I�:ͯ���,/�gf'�&/,Na��IzJ�إG��;�[�9�s�϶����`�sQ	EuL�zX��62?�h�r�<��-��'�����}�n����c=���?0[۶]8`���g���,�e��_�u�7�ؙӼ{k���fk�p����g��oB�y���8��'��\�1SL@%Ka-ЙX3��mι-D��q�p��(����e{��
��\G�j�N����E6n��Q���'Dy����j�U�p��~���ml�����I���^8z�$P�(Xpj�P/불xe �c�T-"z�5��x�O*9E��C�N:��N�/0y���S7��ZN���C��ˍ��A6֬�K�]�$r��jCEQ���Qq��J�E����#5a�N��С���K��0�_m�y�sW��}��9�u�}��M�x���}`��&z�n�~���i��ѓ�znJ�-O� ��m��@�.�y/ ����0d.���i��b��:�B�Ƙ(���d�w��n���N��Ծ��M�ѿ
�����q��]�v�.�\��{ʦ�j��[p��{@����ռB'�#��@������X�jП'��H?ƕj-dY���<��UcT�
��s'�!�3�#��,�G���3"��u��\�~X��e���6�wj�n����E?U�A�CPհ+����#o�Jw3��[�q��j��gy՗��s�F͛�c<�k6g ����|���kα�Б�8�$�o�g<uBԜ�8�y�����zF��-//��S�p1�'��c���)�of�>:.x����u��}qt}�&D����.h%�����{5���m�o���uϓ�������-�{>��?sX\X��(���忛���|�[�C���{���m�o�^��i\��>�9m��tr��/���I����>����̱��<�[���6J&$�7�����K�����[��Q��CA ��Z�}M�
+�D���bm'IEI����U�T7*�b�%J~O���\�;�K�s��%й��8�/D��j�!e@>�h:��:T��)_e����x+�cK�h�DUⶹ��6X��Iƽ�}�]�B	f��@ŏ�W6di�'�B�bo�'X�z�86(�I�0i�p�����x�v����9�p�ݼ��+�kW/٩ǵ��k ����'o�/�o���G��7��m�_��-:����'����±�E��W��� ��d��r{uP�MB��!��ww��#����IeV'�˗��w��ٮ�+��۹sgl�����ol���59�>�<�x�Ѽ�m���`��JVr��r�u4�����H`YD+�m�Z}	�|R�N"�C"�� 1�=Oؾ��w�Ҿc��z_�lH|-�&�����l���] ��q�S�]CĔPɑ���?��q�)y!4Mɂ*]�����Z�bF����i(����t(_�'�<��"O�M�l���e�B.�ٞ74W�f=?g�~%�|☝={R?��s����T(c=}��so��K�Ay�
D�+M���>)i�#Q�U�&�n���~<8=���{�s��`e�W)�;�[��ӿ���L��Z�E/�)�pna)����c���^����/C3��C���`���ZC�2[�ԑ��A8���ͻ�8�Jq��ϭ��?�sKI�F1��b�'�|�B���QIE.�e��:�Z:��m��t�vs��,�[޹u	.��P=�BK���P,�j&]��F(y��$��;�08N��"o�3�p!ᕥ�𙯾{_]t�1����X��nܢ�Y-�ƾ�����;���G�m��J�	:޽ԛV����lw�\��W.b2���Y>���ٱ�6�ʯ����~�顽|�^�)���g������R/Md.rȤR�O�S��1bȬ(TTB
%"�v�4��T����l��r�][8�tn��.��+���W�O�޶;�.�ʅSv�첝>�h�Xl�Ç7o������'��1ǰ�❥]����b�4օ�������6p*'��Q(K����95a�X)Q�N�����D�Q�jQ�)���$�[�u����^z��[�z]5	�� ׏^���4�b�ך�6	%q|z�_*{�ً��׋hFM�|�m�T<);��'���R7N`�ʸx��	�A��옟p��8�ُr"f߼T�����Y;w��]�~پ����K|���M��>.��l�� ���s������:�N�D�-��!�R4(2����{��H�V �:�D����9įY��2'�@��4�����\�H8�rN����Y��ft�N��_t��-���={��6�6�p2gpN�s��bl�je[�
%o�+=��0V
�k!�t�(�e�7���έ��䲘@��n��u\�WQ�G�>�(����ӘgK�s~��9���!A�>
��:p�QQ�Q���Z�FU�:u:��c\�ؕDAh���!%Vq�:N���7�Y�V]fDfr�������s
��������@YP��t��!w
��Ҽ�#�z�]�t�Μ>����[��������s���׶�N�ХsBi�q��;uY��8���G<���^�2?���u��`���bX@����¹��t���Z>���4cgϝ��7V��[={|�4�v�Ԓ;���?�9�:�9?�~����B���㨎v���##%��^��،SCXID>������8�]I����>�r�t��M=|�<�nxW���C�P���wF�=�/H�2H}��~��I&C�Ib9�G �qjt,z2��aP�T����F��7�K�tLA�g�;E���r�#;�*�@'�+�a�!/p�N+���l./�f���8�l�&_�qٗp���֊}q��ݸq�Ο?iǱn�*>N���xA}����A���ql%/l��(Y��"���JAn�]�o߽��<���#�������K{�f�(�7����E�~��ϭ�����'lf�śN��� ��@2P�J'�����F�"I���@[{f��h�VY7�A�	���ZG��Q�i���ž�8 r�*
(����|���;� ��vҢ��,�����c[���w(�-e�����.��\-�~o~�^�2,��Ug�E��Z���y8�<��#�]>#�aۛ�����+�=;�+�gOۥ��̩�pv��o؅�����Ƃ�˽gv��'���;�X����7�y��B_���g�6��@!�����]H�b�r+yGે�O"y�T���>��w�n@�M��޵��v��I�u��nx�'�8f���۫�۠����{�jכ���U��s� y@���D�$����a$�݆Jz�"Gܵ����;��&�NB89-g����IH'��r���.���Hs�
h�[��B�2�&��c�'GjF?S]��E�C�[?�|�בfuʒ���.{�5���_(Uj(�mVm{��,��9��[��H�H�6�O'��
��<�z�y�q���'EH���v\)�zIOHF����2f�f��	\L�^��'��Ԕ�==k�/��]�r�Ν9asӺA1!�!�i�����1���� ��d��X�`XQS=���~#�;�Mxn����>��f��;m�ۦ��~���}��=���{����on�����c�����+v�kv�����h�sw�ec6�8�+]\�z��9 jۣ�<,�h}H�$���i����F�'z˲H�ʹ��#e�:����1��:�a��hmi�)r(Y9���!W<��
@�lYI�q�H�r����Ѭ��x�B��̜����8�y�R�����[S�'_$	��(��#B����ꖝ�Sw~E5�g@I0�ʹ��\:�Nv��׵���%�W��3X4���Kg���y�p���%��C��d|��ً5���5ۧ���K[[�"�Ǳ�4�jY�R>fJ�$E�x�+$��G}H���;�뎬�Ғ���a���aQ�ۆ�cǏ���s�v��E�u�w��ڙ��mn���2,�f�k{���=z�ʞa�}��}������i4�S�Ԩ�U���'���Z�R~��,�����^�F���홵]B�������m�s��-��Иb�kXf�e��\�u\+�| �\��,�yl�dE����*�r?2@��l�} ��0"_�`XQ�Zl�	�K5�ZT�a����f��OB������8Ѵ����.�T$ժ�)��m�o�o=?$B��]�&B��J��=��O�x��㥄�87j!�Η�C*������ޔ�?3�x�]�|��ܼ��jE����a%ƒ�?r q�G:����+l��8u�\�֠���������u�<�
�j�ٺC��[�q���X���{�<za���p���x�a���f�P9~|�.]<�>q�;��S�Y�ߓ�qmg{�cKö�4���qx�Ɣk�"^".�n#Q�)�w5r:��H1^��,HPG�4��\���$f�H�'"/�i��.� �Xg�Z���˳2m�<����i��n�H]�l<`ynU]����h`��7��w�;8���ϭ�+�=.���'�+Ye�X1�N�����ܜ`}1d㒣�`��wฺ�Lgϓ�?[�����A
>������!�Y��$�Iv�3ā���W��R�O%��Ea���2d�
�g䗁R@y.�����<�g�&a*�\�ܱ��Xe��[^��J4'p�[,#pl�ٷ_ݴ?}s۾�q����jʱ��^�����3��_���߷�O^�ʚ?���*��-�,�MAI�
�A��ݽ?�9�Ʈ^}�~�B�,��-����.g�?x��D=��� c�_S��_ǉc�V.�����a����}��9�|�F�_ln�=�n?������{�ӏ��ŋ7rz�V�Y� �6A�\��y�h�p}2u\���_���,Ĉl�!������Iع��S��εm]��cMeH�G@mC���P�{��:6D �'��cN���Q빮̏�#}�@�<!�9�)6P�r��ԏ#��A6�<��vY.��1�!�
j�B�#�^�W�8Ι�e�]��qK6FB�����w�*a��\$�u���d�9Ψ��<�W�?D����k�vīP,��r
Ik �y���9Q�%s�n2d��i�϶������)���Ҳ�\ƹ�����nia��\ߴ��[}�o}��p��ߣ��G��qm��t�Y�k����b/�"��&J� �R�%x��F�$؄6b>��i�(8l���Xc�s��%;~�}&�v��b�sK63=g�?hkk[ￕ����gȦ9We?~)���8�x7�eg��iv���O���"ZfP���ܩ��o�y����,^a���8�hw}���F(�����7�s7	V]U��B?��������[N����f����^7_���NAq�x5p��dSDD\6
��(T]�!�=hqaN���s��ˣ)LM�PNwA�s�h:�a(��:���%}eM��!�Pں���tl�G`��.L�PF�@C��Q�ԣ���@pn�2ktY��Bt�Ȗ���ʉƖ�2 ����^�E��0:(	�epR�Ur�Z����U�W�`�7���8�P{�/����4����)�qE�;�3S���4gW/��c{������r^wmٯm\��}�e�����C���������(�ѹ����}B#��[| g'קA�7T�@F! _�X/&��1ߴ��H R&������qnm������wp���SR�O���[plo�+��?lz���=}��~����o���?=��O_�:N&8��O�fpQ��!�e�]	�)݅�OBQ:}+Ԡ��z!ѕ�k�$nl��sq_�7��a҄r�4����(��0B1@'-.x#d���ǝ[�늓�q+�z}��j�?G�f}���-�}��@%�n���Cխ	�6��x��/��m�Xw@�_�Q���R�m��xHP7�#��j"��5@��t|lcI	D���ڊ�B��\�Y�?��
33�z�ii�-�O�4�f���f�8������mw�g|��&���]�P�D8���6�T�<J�G疱�de�ݎ �:� .�%e�4�ܢ�>�'����ޭ��F�y8�ǖ��.�Cw�h���ֲ��5��붶�![�Gv�7��t�r8|��FX���VL�1�{E"���\����}�fV���AϺ3��eN#�s	c�w⑖̎�
�*B�����I��47����\�R ��%�f�AY��S6]���ؤ�A�Q�kB.
��{8��
/�d�@^5�q(A�(��u�~��������|��ǿ���:�MR%L�|*ǐ$)�GvIFb�ZtT�eI�����"r��1�5u�򠸮p�ҹ�tI�Ptj�0Tq �U3�AZw�5�I�'$�)�irՓ.�=���������2�}28y)�hI���� ��d�*Dzϟ�]����_~qC_�б=�v�x�~�~������'���ܳ{�>�woֱxr���eZ+�]8��!�<d���U'��\�8���6�8�T��P�6Mp�0g�+�2c�x�����'}o]��ի�t�����k�s뺝>}R����hv��������o�o��ow���ݵǏ������W��ĉ��õ�4���g�o�#�<���F�B{p�H;I9'g˹����<-�(�dȬ�Z��p]?RaD��������i�R�A���?$qtT��dۭ���"������ô/�oSg8���������\�(@+ �.����')é�Q�U�~�m���\��s�s)�k�U �@�#עcKX���5:LQ���Ғ��/��..�!c�� ��������J�?'������Z�(I�0��r��2VQ����� ���C���Z�6��z:??o�'�mq�w���/���������|�����ּ}�*�wp��~�����u����>.qqΙ��"?�vDWJ�k]dU���� �Y����h�� �w�[M�!!�,�+D`�QV�4��Ö�#W���Ϛ��V>�)y���R�.eѹ���12�������>q���2�($r�J?P��cL�:�[�:�|�pa>���_��w[�䏅��\v��� ��;UT*2�1W��ˠ�9T(�)_Nhv�;�R���Qw\�8��ҹ�[r���u9����Ae�dtߝxp����t���v�܋�S7<;�~��H"";F�4z��b���i� ��ωpl����M�����n��_ݴ��/��3'l�!9;����}��8t�������`�z�->�@�-Ѱߥ��94���/r����r��Ӽ%OM ղeF���X�|�E,�EϦ� s�fgv�ܹ�rl����݆c{��Y�@ଢ�~����'����h�/z���'px��-��-߻�wH�+�O<��M]�)�~�<a0����y#�a�G{�rK��-��]2��"	&��&�S����PtK��Iv6r����֏�?���Ǵ���� ���C��&�pߏ"��e(o� ��X�.˸���#�Z �
K�'_��'���Z�7t�ӹ��H�(�op�x!��n����|��F��`^\\��8o���{}cӶ���<�Y�ӟ<��`��<���N�-0�k��=%�Gui�v>S5y��a���̔��M����ҹ-����w��&���]{�v�-��?s��;`�.w�y�����wnio���;��I~�I'�Щ���"�ǱQ��6ȹ��{͗�7�9���b�KK���x*;d���ہέ7�٪�@��έ�k�s�P�!�������d��?��|��(D�6�[�F=�����v��wܹ�/���N��QH�K:��/m�V,�wS�,f�/,Ȏ9��k�i��Awn	�s9��2�iD���jKM��O� '�)����SO:��Ȯ�yCB��P�.y*u\Xd���W��wh�غs;9B1烈�0�{;[�U��ޙ�_�˟��/oڙs'm'e�U,k�����[����~��=z�W�s63g)���m
nG؆Μ�I](�;��w!�3�@:��.�!ƞ�QȫmO{���,��8$��Ol;��mc�x6�u���_�����M;w�-�3tT��nn�۳g�����ɇc��={���f�ќZ4i^ �)L�7NfZAs�m��~z���L��a�A	Q �EL{v��JȦ��ۦb ���h���E���d�v�}JH�� C}w�nfG�{�|9�{��U�am�����iCu?��aگyz� >�XZQ�����U��3�jc(��</9*�:�0���A��$n_0��rFQ�3ض͍5{��֢M���;cssszU�I�u~�E�S���;��X�����~;�?c�(��V4F'YNVۄk[�����8��t���Bf�"	�������6�wu��P..�zt����;�<W��-��m���X�as��c���?��{���GBh[�7���η���P�I��[��vu��C���q`9�I�?�{�3Kھ���y��9�=灜Q�����#��"��C`i;(��<�ե�sn�ah�(o9�=�2\� ���`��y\�O&��Dp�a��j��(��T����̧�!O�$�D�� 5/�>������[���ڒ�d3B�С�u���=��tp�FC|�!�f��<'N���E8�gϝ�ޅ咷�1�'������ྴ�/�b�俘�ctlsi�N��n���?��X�����2I�(��v>*�4�p_�X���nd�|�B�9�0����x������-M��?mׯ]�V\8F_���aG���|K����ӏ��݇���k-�\@�cI�h�cu���2S8����4�t�x���أ&`���� k�f��&X�����1�������Lp7��#�򒰣�#P9�M��Q���!`��nF����x�Q-b��R8"X��`{�VW7������3\\?���>�����;�o��_053aK�f��������[��Q�j\�p�����yzf�D���:�~����J�����b���w޼~g�=�_~y���3�.���:��l��"�k��*�������6??-��~�5�>��]R���G�5[�� ����y5�)������n/�#���Lc-d����i�<�M;Fs�H�.��%=A*εݳjvf��n:��ԥ;��w[�]��+>�t�����^$t�+ ���>O�B���1��_a�>ۧC��wn�ǅ���r5p��� ����2�
{�e�!�gVg�H�+P��3�&��Z�3X8�5Q6l�;ش���X��}��M�}���9sW��:a\+_�^�����������'Z@v���wݥ��#Hg��'Z�}8V�⊲��9�%�e�(�}X��|�X>C[��6����8�8����SS[��hv����tǾ���]��b'���,d�K�%⧟^�_�v���ן��>׿�Q>�>;7/����:)¶9�����W����z��R����]B)wC��#
ty||\t�\�{245]����b��dU�q�/j�>%�mpt��WD��Η�Ȯe	�Vّ��F��l�c�P��~P�]�t�yϰK��u�J�o%Ev��`9��
z����x/p�q�����t�5�k\� ����UG�K��c��83�!��æ7!��6m;;{���[����2�s�l�*`��ظ�9!�
n稉+|���4e$��!�mI�a 6���;�0���;��[^,-׏��<2�E\�݆�8gM���_�9�?��ɍ߰��Fݡ�l�Ϻ��{�=~����X��Lw��� �����^�:�6{��ϝ/ }ң)�etgZ}>�A@��	��y��E�12�'�['.���[���TPv_��][�l �O���sKʊA�����\���xq��wnO��/��;\4���"N���k�+��4��0*DFcz���P�K��H�;b����������hbr�>���Ď�;��$SA�!�A$sHuB݈���*���j�5��A���PH.��d����@��k���2u�-R�P$���-�6�-'t��?��=n�|sK?$�|��-�c���[�ص�������=8v���3����6�E�_������+`X��ۧ^�rJӠ�@����(W��7��Cr#T�n?>��*^�����!���Y�����-N�����֭���_؍W1�O����qޮ�؃Go��?�~x`��=�7o����Ş~L�\b�Z,О�`� M�-����LwnS�$m�O�\Ć������bw{8�*�����E<Y(K�Ť[�1=D�=�ةnA��XH����PɯB!�O��𺝵(��&���G������q<Au?�z�Xh�Î=x��.q�R�mf�B�ݴ���B_�Wbު������3k""��Q�̗i�g9�G���>1����(���	9jN�"�����>k���.���˷)����ck�I!F�A�p��]_/&��q����N+��Ju��*�����h��+g��ζR~���cpn���"�x}R>j��h���-��ځ�u�o��	f��q΃C����Ѿ����<��1�2
n�C�uF��0���`���ל)*��zӷ"q>#M�C�g��O}�3J��G���C3�G#�I.�UV�y�1��X�r����I���2��&$��(���խz[�a;�G�
AD�yn�^䅲�G�8�@t�?������������yW���s�@":�4�;����Vlz��I�Th*��s�4 ��dcH9P��1��Գ�tNy��2W�k�i��:��畄�N��
�L�Z�OrX@|�A.�2��L��Jl]��l�&��g_���Zq�A>�TO	��눖�MɃ>rlA�;��hjbW�fK�3v��9�󟿴[7�ڙ�'l~��W_ÿڴ����s�+�綺ʿם�;��?۔]b����(�n�v�X�`����}i�s�)a��͜���|�uPq�6c��=[>k�?i����޹sپ���H��98��\�cK����u������ݳ{���۷�6�	�w�����,��7#���o�y�-}��!��)�q���xKnH�	��E��>��,�\�0�3��
��PF��yX��k�`^7�Ο��{��ۡD9��������K�����j�M�X�u�Z��c-Ka�j�N��4�/e�B��C��X��V��S�=B6��Q�#@�#� 	!D%���<�5�Y1�1_˼���B��S����Ԅ �c?a=����K$@���sIt�����)9�rVw6 Q>�Z�3��<�g�A�;�8o�.����5ۄ��?D���.�1,H7<}�_���.��񉷏�r����������s�|�q~湄�^��7U�O�gscC�������-/�[�_��^��f�X���<��:[r�yN�@])���}څ�mMq�'r|R��1�u��%A�WB��@�����dg��i��u����K���׳:���h���2���ԗ\�1`F��;n��U}�2��2�C�q�A0�sUs��)uR�W�s����(k>��f)e��眅�3u����� ����"Nt"���	*#�$O �7�Z:�P��t�@��K�1�$�i�K�c�#бu�V $�L�y�I;�4>��ppU�rn�d�� d]�!-g9�q����@iesP4 A��*�H���ʩ�g�X�W-��,�*��ơr������Oڭ[W�U����zƔpwg�޼ݲ_��zb?��О=�?k�L��L-F���z2��c��Ӹ��B�8Lg�
tsѳ�P��Z�<=C�N���kR�+�m�â����N�?ٿ��ݼy�.]:oǏל��A޾۴�O��Ow_�O��/�<�/�ɱ�][:��`�B��BR �Ǉ� �-̳��RR����mϒ�A{�� ����n��V��%�y�C���>���<m������C�k��Tu�O��"7�.A������"�v$�OD��M����m�#u�sT����bSY�c�c�3��QM{>��[1 ����a�����e�ӡg%�أE(g�Z���y<�7M���BG9�t\'�q�ݱ�o:��t�����%��_�O��տLB��B��/���(�|
�j .���ϳ8�h��^����L�yj!b����%��T:F��1p�����,��������ĿH��f&�owrp&�]k� xcmS�`�o"�GHD�v[�s�k�~���v�B���X"�<A>6�6A^�$�n���Q�q��:�"�rvy�U#m�����B'֗��!�a����~/0.�Aˡ�.y�����&f��A�:чaY�C�O""�>����_�GY��|K���Stn����m���?�q"H� *!���eXN����r��R�'��V�D��yǜ�S���y�P����Z:�,����-\��QY-p���id���.�e�2%�'��u�g=2Q�BvI���h��
��N���������;��oe��.p�v�p�����O
n޸����3�z}��ƾ���~O���'���q��mt�&u� p�1.�'⺢���b˯�X�ή�J3׻�n��-@���E#�sf����.�X��6�5���=;w��^{��֭�v��9;�����U�~u�������g�ؾ|�^����A���-vǟoc��{��Aq�0�典�pt����OÓv*|8?�S�	rS�dfX���hu���X�$���������}�(�yoՈ��ͺu����V�aa��͉:-�Qa\a�3Y>�� ��Wo�.�@ %(���ҝ���ʻDd�E��ĵ⍽RW_�������j0���!_��.�U�#���򇴌k�Ź�wnwv��B�ٹ98u3z��k:O��X��fy�w� ��m[}���VW����W�n���]��2Er��p���.;A��x7覓��^S��K�ZG�Qwt��62��<����¹]�s�׃M�ϼ�������<�۷��f��6��_����2�{��pA�F�ى��{��v��v��뺌�4����l��'�rncn�pSkD��M�֝ۘ���so�QVqL���(/�I�ǻ�)L�F��gn�s:<�IPW�v��*�����>R��#�y�J :@ſ(V�Yl�y���~h޹�G�#�NQǉ��&�T:,猨��]S'�g�����>*�ZU{���e%��C��<(�"�|&Tj�n�]�'e�@a>'�R'wp��o'N��ի�ڵKv�+�+}̈��{�|��?xiw�>���ַ��s9Y����x���S^څή����<(��^>D[��~�W�Q~="�z�7����n!o���'���E�����+rl/\8g�Ǐñ��qL��}�j��¡�ᇇ��'��oF��	d�}���
{�D=C.�~rp;�� �N����E�A�7"ys6�1ய��������K�i�t},���8��h�ߎˠ�q��u���=`�����bX���H"O?%���KiG��0ւ�DWF��6��7�C�1�M�y��2��~u)r2�ԝ�]���M}�rI\��p��g��mړ�����/�<���ǿ|Ɣ5�'=�O���œX�V����X�p.��cv�7mN�tGN���;�t0���M]*=e�1�: Z��*n���K���h?���<�IӺ���;{��=}��޿G����������������"���y���@�N C:����PW�P.��������(���z�'8�F�=�V4�M�v��$�n:��n~�e~7� U�TW?��*M]�c���k�c	���z�
a�$y��I���y'�2(���q��(g��d'�'����-a�F���P/Y�AY�s�4KxU����;������v."C�R��/�A�@&����=-�eZ\�V���k�Q_	'n��E�q@6
�c�Gx�2��ى�y����u��e�g9��6�_o؏?=�����~Ϟb��W�|_��Vjqk&���>z_�6��_Pv�kSƉԗY��"/vւ����hj�3ڂ�ӱ���@�@�-����W_^�o��c+�/�
��?:���g����/���o?����nl�b���ƾr}CO5]H�e��)g��"~�$���Y$�$ �۽�|"�-[a�����(I��n������F��,<�*�H�_:f[��P?{д7���'
eQo}�ש_'�s���������%��]�m}(T�C��[�[տF������(ݽ.u��h��]���h�JI��r���\"���q/`�'�,���5#5/2h?��N��ܰ��[�������3�2�9`~v4��i�K:y�����X׸�m��� dS.�{$�s��9���w���ד�O2u�*���2�ĝ/�"N1��ycu�Gt�7ӻ���f�g�եl��;;S����u���on�-_�y��a�C�D>��[5ȶsE��$�l����?2r>x󃨎��JU�x9B��@��ێa��[�	����c�e��y��K�Mwn�ا����~�;���dZ�����A��GEH�^qG6��zu&�[c�H��HU�`�ئ�y�Ch����3y�V�D9��@9"*C�q�@�s��eqe����^P�Al�P:�E(o�WA%��좋��G%5��^��j��/�F
�����I
������%��M��s'q�z�.�;GwI_]����z�nw�>����=��G�{\���b �}�;��N�'�غ�ʱ%/��\��1�.�2�)��.�,�8���w�bq�G��l��<��Oٍ�����v��i���3���E�v��?xmwyf��?�g�������s�N.(�[P<�������!E�wpu5���y���^�k�8��K�k�6QF<��KaP�6_����F���R�F��ق�"�x[�Nm�F�<5��>Xw����v+�� 7R?����}��<d��-]�
�}�CO����"E���G:�61�u�$���I����(����W�����g�+��\���������i������sv��������q1߁���a�M�o���$}M�q#��m��e�tˆ�G�H�_v�	��c�I�a�$���?ֹw���W���q�y �:���0c��.���q.��z>c���'xN���|6o��Y���^W���� �y��$�1���X��z7�E�9����Hym�cS?�$c^c��2tR�XJ9D�-P��G!��j0F��}��X�eڣ�&�&7�����*p��BOm�����m�i\�l�N�p4F)+H��j�ɦ�������1��sF��`�o�����'k���_��*_6��W�3�_r�ݤ�����=��$ڇ�&�D���3����˫���hȞ��5i>���w�ݙ�������<�d簘]�|A�{��-.̃�*�W�{���������}����ܿ�M�0xCo�#�$��0�����a�'9��c�PcT/�1��Zs?7:̼�YѸtA�r�����ī㐟yU*@NE�����|��W�T�.QG����@�
)ҟ���TA:��5
y|��W�(y��jB��o63�x�i������P;�����y�@R>ڶ�φr�<�&��F�\�x�+H�=J���k�N�pp'��ML̡�m����o����Z��x�ѽ���������]<����M���ھ��]�xڦ'�lkcM��kau�7Z��U��t5��;�ُ�?��&�Q����y8���X�x�fJ:���k�����={�Ҷ��e+N=�9���Y�e��I8����W�0�g՗8Ǥݥ�A8K�b�#�;2B����q\�H�FK�K�:]�8��,J򝗶�%� �j6�`_�aNL]��_���Տn��ɼTj<	�D�I^Vၨ��<��.�G�<������&Q��L����6dI'Ȑ,I�^�BY���_�Q/�Sĩ'?g���<��n@��2���-�_�C�dP?�X�I��*"��`M&��r#}\'�q��<F���a�ĕ8������W�'���ڕ���o�ح�����Ӷ07/�յ{�xN�����'����1M��ջ�io���Qߨ��	j����q�p�\�BŢ�c!C��Jb������D�HbC}_\�ֳVׯ]�/n]�;��څsgl��h�����7o��ؾ�~j�ù���S{������w���I�J��6�l"����\�&���Gڋ�a���.�}��4�lN@���HQ�m6��/�T� <��_$y�����%��H�z����P��ќ(�{��&�k��v�-�C�k��@~���Q|���cyKvU�h��z%�}�Q����`,F!
P��]���u��P}f8����o�r�@���(��/��d)��2&=#��Tr ���A͚VG-'�Qb�/�Ր�R�r	p�A��_�y�D.�:�;��td�kz�[s�������?���������gp\�`��EaksUi��;�����F�N�����NUO��s�����lق:�N$ڝسݽ8��� �?0;��-.��|�;���nm�b}ߵ��u�E��7����R�=��|a�a�n�NR�ˋ��ODv��l}�2��$�v�y�ě.<G��Rx�����?˸�Λ�k��u9���M��O~ԓ)��!M�!�)��|-�ҿw��JhS7U���
��c��y��lG�K?4�eu��E��׏�7��5	�`i��%���+_��߭olAh<sY)�>
�1�Z��)ņ8a�9��b�<����#Nh.`N�O��/έ���e������:p�0�sट����_��R+b�<'nĥ�d��6e�De�c~��z`O�֤��<�Nm����.�y�\l�M�>�-�N������*�Mpm��ܞ�9��v����m��o���++X��%å"���O�o���髬�Y�i@����$uT@k��^��^��X�4K��{u�jD��@���6��ӎ�3��U�a8��{�_���][>>kWV��?��K���[��K|�[�c�o�����Ǿ�g���Ğ?{�j𮭿��0M;��K[�4 �c�}%\}���~С\�,a}���\₃4�Y���`��$$�q20)��'����Πm2���ц����go\+�q�1sf��DA����:���$C����~����t��oTN�>6�S>yz(���P��E�R7t��y�*$q0����HP��v��{�샏U�%(�,�@C��s2��f1��~6�]ȋ:]h��( ?e @��]�G�l��O�>o�Rs#)��X�1�ǔ;��pq�� �EVC�n�?��P��'L�x���8��?*���_�3��v�N�X�c8����j�(�G�3ǥf}ݟ���u���M��h#�M�B��Q��g2d��L�i�� �?�bi�y�M�"���"�;�(?���.m����m����۷pp7d�����$����3Ϸ`�A��JRU(h��:&���V��U���>W�5����>isLy���n$&(� ?���G�g|�]��u,���~G��S^�J�t����.%x�,�����qE�����gn���Fl��)���<��28(^,^�-�f�$n���)��'֣jC�!����:����u� H'H.I*�2���<�3#�UB�se]a"�̮)�z������#���(Eٞ�݅imҏMi�,lW���C���ܦÏ8��yDH�`��k�r\���_�ѱ��`��4���	;u�~<�;�ϟ�Ǐ�+������ߵ�/��ѣ7�4��lc��$`Bb�$�� ������d��)T���N*NB(�> 4���r��}f�eG��k=�{r�vvݱ���D��=!{ή^�`�.���Kp�'�������>]�{�^��w���{�a�5؀�y�wJ��]$~g��s��Nqn�˅'��|����Jv�����IN�]���N֫x`��[O`Zl�B#C�-���{��^Th�
,`�
�IQ2
�oe�w��;��Si��y>ꄇD�����n�O�TDŁ]cf�N�3�qjj�¸��u�~�&�$d��X������0j5%��lh ������6���$ C�ԏ��Jd�ᎈ糹ҮBdw���z��ǡ5Ak�:�5O��/�� ~�4�5p�޾��z���?x��p��o�m����n0���\�|�n޼`ׯ]��	|M���=�w�����x���p��ԝ3>�e�b�6n�u�yU�x��\�m��z�j�����^���8�m4>���⌝?�<�p�Ē����$��;}Sf�MN��O���9�
����k� 9�ui���p �d �k�k��N�Ѓ<��������v��\3���D/���J�/�	����!T���_K��e)��<Q4I�O<n�e�%�������,��L�S7D<���
@���V?S6c9�}�s���hP�6�''��d`V.h|i5�gH���U:�o���u��Ņ;sfY�{��98|s�
e_̶6�����=z���o�޽��^�h���FuUF�6�~*�r]U�KGC�%�P�|����û��|Y�,�F�ù���m\��صk�'�!���|��g�k����&��g�Ï�px���1��<컨g���>����d�>Ǐ����{��t�(��F8�#>Ӷ���s^������VN/nF�ʜT��!tm�_�,O �A��p<c�bi�mBP���.�����y-#?�@Ԫ�~/|���ϵm"T�c���S�vΏ>:���郺�����@ԓ��C��nϯ�a09.�f�����6e����"�H�?�>�-���r��+��y3��)sT� t��s�iZhNdH�qͻ�|M���l��ԍ�W�W���W�/ޱƭml��4��:ߒs��]�z�n޺hW���S��l~����d���?���$��T�
��)/ FA�vU��ѣ ����AN��6�w��{�n�����O_ٻ�-�Ĺëy0?�~y^煳8?�N���c�;�s� ���8'���fO����Ř%�r�^�xUƹ��EfŐ��
��9�(њ��8��GG]��8Hv���r1Q�#������\FA������q��QȌ�r#z^���>9��5����:�.GE��u�f��"�<@�~u�1I����"o������ˋza�������p���X:�fkk;���{8v��ٓ7pn���+�#�"!�x�S�ſ,���V��Dc;$sV�K����s�BZ�|��	�U��ם���/���_�rQ?$[�!f�њ��]=����k����z7$E�/��������z�m���l:�H!^G�ԝ �N�6�Xx�v%/�$���y�C\�rlh+�,�:v9��84�:ݼ�?�G}�&�j�3��!�Կ_4��v(o۸�A����>�ޏ�O����9�6�$ЎaK�3p�Ҏ��:B�z�z��ä5�Z�%M�O��<|o���y�aO���_~}f��{a/_���:.����f���,�I�M+vi匝8���:���:�[�-���I��jD���GG��C��w[�#�=���ӧ/��c��=�|3����?;3���Ο��{Z7>���[:���{b��7���q?�~04�:���l����ڭٚ�:}�ZҬ) ��'�Գ֗�D�ח߃�Q�I݂s�;����F�x�2<,X�D�n�b@���N"���.��3A�(�5��6vb�ܨ׭�aN��i��0@zʬ��!��ZQw
�_������3g�گc��w��f/��)�����v��c{�����r�=\1=��D�Y��5&aW�]�q �6uf�0���"��λ-|���}mbb[/|�,�v:�wٞ={
W�s_��k�����+���#���v��3{��w|��|�C'>v��=���q0��`Vɦ|wBE��%�>�c�wǳ<DH<�&��;B�?2���l� ��0��Ȓ���Q>
(�9i�9��"�����ǧe�8�1�&�b7����>i�_~����'}&�><6t�����&��`]Գ��� >ۯ��8uT�*m�AQ>�l�%�.��<&U��~긢.�sc:��{Ac��<WR�'��n�ܵ@zҶ���������v�קv��k{Go�' �5��V^�۷���[���S6��ro�����;l\��"��Bt ����N�r:4�J��#s�2(X�a���-����G����7��݆~D��h����ų�r霝<q��it��Z����)�_'���3���n��P��!��E��Iߢ�>�����<*$�̩��P*��F���)^�oB�J��:����e<�Y��`�R)�=��~Z�Tl\t�bFi;����c�;����=��ReX���4�?���c�*=cg�����{Y^����������;9���}��/;`r�,�9��]�ފ��x��	;�*���a\E�Sϡ�ߵf�4Wx��?��5L�������Kv��e����%9�����枽|�i�r�翰���|"��y�Ý���`ЩwG��d4!L���O��{8d::�~ޞ���X���'��tdG�ބ�i��}ng�Q�%����U���4N��]R͆Z���B�+�&O�c0d�?"J�b��7 L:��xj�Ǡ}bG�v�Lm��a�(%y>����?�:�\:tl�C�t@��̔�:�@��R=�~orp]��ξ��A�����}{�:�/W���W�˽������a��gf������3v��%�r弝8� ��ğ�6�H��>��
���pn6��Z8��)6"��S\_}��v՞��}.��ex��W�3�M�5�pᔝ\^ҹsw��⿶�y|��[�>�e��)�D�a��CY���|Np�`J'ƓXF��#�@���J���rxL��,��6��ϡ"R�k��GiP'�[�Vu�HL��L��c�6&9@Y�	���P�CJ�������W�\dv�`���ꝋ'� ���]ۋ��ٳgʯCiZ>\��n<��_ۦ[���<ͷ(���/���o#`�n���oMVX�嗸�!�P�$T�����-��޳S'�������_�wn��S�X���>s���=z������jo��o\L��lĻ��;m����;���/J?Hi�B�i�Hff��?�Ă�vt���˓ 6':����N��y�t��[���>�c�)pL�?G���x�D���SC�@�	�"�?1��NJ�^�F�� u������3BsS�:��&�Ǽ��qǻ�~�U��^T�q\��3]]�N`������k�.�Ւ:u�r��	˼d�������T�WeNc-��� ������t�����{�n]�A�<,Crd��^�v!�ޞ��e�3��lk�o�Y��Mم���I7!=��d�!�����t;� ��rG[):�)��Y�g�66������#�w��~T����o.�֟81k�.׻�/\8ks�M�ֺm�����u=��G���"6���E��"�C���7D��9�]�eu.�1Ѹ0��ԁJT�����}
�ҥ�X^t��I%�C�ș��B� ;�S��T��꠺㬦N"D��u�Dt�*^��>I�E����0M����T�,:*�ID�'&���'�&|߷��;}zY�����ɓ6==c|�����=z��=}���^�<~Uï� 2t璎���\���騆���,���rk}xܦ耫m�&�h�pr���?��c{��9��7CܸjWV���_�^���Ōw0=�Wt/��×���[�ܤc8i������Gc8��Y�L��'�y{H�*� cNLӌ�7ǒoi��Z~E���Y��f扇c�%�x['Y�I�
�-�7�3�F�G�A3Pύ%��>�}{�s�C��|���m���T�u�*�)��@��:%ƕ%���p�a+�ÐD�t��?C�ܱu��<��q�����X����<���u~9!rDHpJ��5��t�t�yO����dq>�xۈ����x�4�SX�qa��koޮ�chp�=~gN��C7�̖�f���e�|�]�z�Ξ�:�\s�{�&�"�$$Լ]��"P>(�F��zPգ�l�k��^�(
x�Џ������ڶ���ѓ�셿5��eй��O�\�����58�����k���
���-�K�Z:�����2��BPڷ �-S8�(�dÈz\}!9g��Z6U.�#]ʓ\ZCbq~�;���HFZ�ȏ2J��")K:��ğ95o䃦.��~ǫ�=��J�k�<�
��<B�&��2^"��ȤJ�?e�yYU����@"'���/]��+�(�90���.'~�瑕�?~(�+�"���%b��q�Õs�#6�[E�gz������; ����� �(������<����e:�{�
e�Ѿ�>����ܼfgϜ�i�ݮ�}{�������?<��p�V׷����
ub����?��cK}d'���.=v	��&'��@�@D�b��� �x��:�yj��V���%[�t�n��w�ۭ����f����~m}ߞ<]��xd����剽y��xzn������'���ɋw�cL�k)�Y4�X���ƋE��O�-�y�#|��q.�����ҙ����򝌼�N��uԨk��?�e��s+�*�0���c}Uk�y��2�_a]�#f4�CmWW��eu���!���1C��@q�V��P$s�����J_~����V���&�쒄r|�y�#c�)���U)�X��d��J��tq}x�����{:�8@!�'�J\6V�+�t�łz��so@�7�3˝�����C����=y���f����2Υ ����T:���<����:q|��$�2�����e����[[G�׍��)��89�y���Ơ.�*�6��JJaF��8'S���~���r�$��9�>G؟?(^X����;~k���׃���9�2[_[��[�{{k�������W7�hcM v�A4_��P�8e�F���!��^�/���p���O���ה����Y����6���jB��{rQ��]�>�K})�OlQ�~Q�E>VE}�}��2G)��nNJ�~�WC��3��CD���IR������{[��o�#�; !E�$�	uU��؀�ơ���� �c�rc�d�G=R��NV���p]3V��7�/T��ن��6�Q���Aί�8&�4\�P�G0x�1��Kv���t�,��manN_������m{�l�?~������0����e^`p"�]@�;XhA�s$=�GbBwr��6G�?�_G�+�|�1�0��i8�+v����+v����foo��Vw�ٳU�w�����#=���=�F� �<��Nf~�Ͼ7&��z�����BΚ�E�;��f�J��Z ��N��=�u�8*�Pٳ���rR�_��#<13d]'�Wぶx�)N��?2?���T�9�G�8�
��ͥ]Cb�.m&��"*W���焚���Oc���_�Oe�&T�W�E�رK��	H�4Cm,S?rMc\L������=�&�/��/�&��@e�r�~PX �l3�A�CF]��ff�q�G�!W�؏�4�~uS���_�ڳ�lu��'���J�S|<���y�\>g�����o�h%�یmG�9.�G�(骠ţx���,�q��QZi V@l09����}�f͞>{������2Ϋy8�gO�+|���%��la�o⹖|ԋ�Qs"5:
�T�d<��s�P k�]�>'�f�c��8��]�,� �8)�Y��EJ�͑�e^M;Ϗ�L�q���K�f�|f�Ef ɩ���o���A�?�?Ρ�w;�@�s��9 �$\��_�sf��8�$��L���"	,0��W&�r�Wq֡׀���z��ܹU��r�:u�s�q�"y(��}3�y��1)�"(����by��d3B9�Z��"��xE��wA�=,N��pzv��y�|��}q���v��2�[��,�J���ݽ���������}]�;�3�|,�:��A�������O���.J�c��,�q��`�@b��S;7ˇ��m��3n��۷3g���[W���v��5�p������nl�c1[��~~�>? �C�_���g:�����ɒ]���Zk����z���v͆��O֟om����t�wUi�Zk���߁�8'�ɬ�����&=�  �!@g��/�H^���S^ m2��w��%�%TU]�A�����民>q(�(nKf$x��hHfjO�?G)�y�e|b4������a+�;�V�#��� ܳ����W��iu��W7��=����pwr_��w7PWqu�/M���b��D�WD�������˓�pG��|�`<@��� Y@~c���_�@u�F2�1t߉��oO8('�.`R�72b�����q0j��l�/�d�|�n ��(���&K���Oaq�l��Uɔ�w-
c��؄�s�5�Oc���0�mY���ү�/c���3�����en[��wq/��J=u�L[��~�M�a�5�dS�n���#O����/:(��Ұ��a�z��f�����<mo邏��G�5Ͼ{<3���Y�8�{�3��c�o#Li"���� "P�2�y�R�΍��1&�%2��}J���h!A�^�(#�	�*A��iewg�<�A(�\gֳ�vr����<:#=���*?��D�I�U$���a��s�ӘjlL�sS�����`�N������Kʅ !Ĵ3����R)K�ĥa
s:Nym�K�B��+���K~����e	��;)�����4�Pn�1@�:|q
w�C�1�I��"v}�щid�'��ΤgOW�W/���496��� ��S��:I/�J?���^7^�3{�?�6{�'|^ˣ�F�0!l�M=ū�R�-D�26���nA	�Ϳ3@�m���xၾk���<����ۇiE<OM��k�xf�ǋ���N�ӟ^�~z�>|��S;[Ў��f�6.fm�jL�%q��w- /���P���K�0#^�GS��w����s��s��Xz13�����U���������������7�����>EQ��H5o@����Ȅ�����G�|#T�5T
�g�}�����"�K�/�?+Z᳕_����7��K^pG��|��'����_I��r�l�@B�-��I���z�Ȭ��2Kk����N"䣗e
p�[�9�ɘ�[ �c7�~�\�(����}�/����,o�8�������@�P�~��܁�A�1�{Gǧ���,]H�S�1v�q��/�Kdrj+��x�A�Ug��2�f���4��uv'�<�o�X�12<�F�܎�H�����������E��ڍ��/Tjz����*�r(�$ت �h�F �7��?��t��M���Z��d�d~C�������w�tv�=���.�#�9=��4�	��k�q(��͔[�$`�*z
1B��B�U�gO|&��Pn����3�z�c�z^k�����($�0AE��
zo������A�*?!SP��_C��`.�L��|�!��xn
L�v�6l����'��A;�����#��;֨`�Bym�:�ˋ#��izj(}�����W�������W.�~?<���w����I�������O����˒R��N�*�y@2 ʭ�(��bb��
�AR��@��)H7`��5;8�k @,.L��Hfm�.��Q�0S�i������ҫ���13�<��v�@�-��<�� ���v���lbw |nO�w��v��Th�,�`ŖC��Ƈ���������}��������3)����R��Bˬ>��eaV�||tAၬ����$�zo�݆W�Բ[)��W�z;��ۄ��/��U-P�}1ﮃ�����i|i�%x6��+C񯜱�a���:��M�WgqGʛ������5i�Ɛ�xӒ��/��Ҁ\�ѹ��wBy�2�Ĭ.k�5 �^�r�vjX�: e��c��#��z�q~��#w�{v�;��cwi~9������Z��3������/���а��!�`嶿�J��舅����Ɛ�trx�It�2>�Fx���!wdf��oUٽ�?�4 �4�#�:����I�Ȍ����x#3��)�Ӡ����,"9)�}��B岻{�O=�ig|��<�C���qݪ/˵LT�(�a"	ŃpA)�b�_�[$���2w;�{�c�_��K�~VD�r�N��e�n���~�	�9BI��p2@M��n$ ��T�l��܉'����̅�@��3Y��V���9x�E8��7g��F�����ʟ�FH�imfh�m��>7�]Љƻ�=<����[*� ���{${fC�d�G�=�yd[�Ѵ��Z�ؔ��
�'�˴�q�޿�Io�mJ���Y��g/��[�?��1�E�"��Ќ�r��@�~?0�pqv��xn�4#H�}�`���NN����^^�t(喓�>��wo>�͵m�l2SmV�7���"�ZY� ��$�3f�j1�;�n\������|K�z�`K��ޫ42�/�v<=z�����I���^����{�u�����JTA�~e*:i��+�,Px���l�J�v,P�kϷ�;e��+i|nz�Ơb_�;1����u��;����+�5�ks�̌Y�1 KQ�|S�$H9�?^w�_MNM��������ۊw�����b4쏳Pz�9N��Q�gz�Q��)�
��"h��L��}L�1������=���w�y��wPX[߱2wy��HiDJ;&�����w���뉀2����0�	���
��|"�X�r�WQ��n���o�7RJ� �R�p�5�>�A���)��D��R�&Ƈ��կ.jL�I���\�����TN?�T�TN&�p�t7��Y�-�B�W�U�	-���0��J��6h�,P��5�/�f��Y�'��n&=�����-��F1�o,DQ�;@��x߂��3�Cǂ���]�eg� +�F�L���N{Û�����k��|o �^���N�����ű*�R�݈;���bZ���GV���+���S��_~H?l����t��6j�e�WGfF�'@:�^";nլ-DT��p��Vh�i_�쐬?��0C���k\�~_<�͹�i	c��{}n���M��=O>mK�_K�ґ���A��Qn���D������y)�^GW�ѴE�u�nAC(ܺȃ$s�|��(��}7��z`�	E���477���zӘp|���|��i���!�C8~�b>��<�:��\⮾j���<��T�9\��eP֥(Kq~t`�	Q�c�C��Bτ��	[�e�U6�n���iD�u��+�G�MT�A������Q��X��^ԣc�ivn6=x����������H������������5����9��=a��ٱ�z�eLJ(Q���T(<>#�Cm��-)d������CjC}����>�`�޼Oo�J;��������'3��R�؉fyi6HB��>��%�o+� ��(�"	vp�G��l�����CnBb!3H%���Ǟ�׽��K����'|PM!Ա,�=�W��<Q4<�5ہ�_Xdu�5���U��]�����V�8,���#�C���Uw��g�(�;� R�S3�!�#}'!p�U�� W0��В_F;
�}�,��p�e���[��(AC�OoB5<��7��8�|2u�D�w@���EX�D��LS�U�t"�eA����1ڀ��P�x�k{d;Ph�܅�W#4�>2�r{su*�����Tz �vya>�LM�a���u�r{p�'�����is{GO����^	*��@��"p������jw{���y%��CI�m;n1P=xG:,EH��^k;=9��e&=x�'l	���)�}�B��]����q}/���4R�zZ��G�R���kɐ^���U�zpH zh���v��%����\��\�O�ɒ�v@��(O-��O��ibl8�ʐx| q���O�}�)��bK�H�!wMo�+���DA��_[�;!x��+�wW��V^�t�<�loæg:����ࢢ��	�O�w��ftU�O[dm��/���H�������g�j��m����K`��ҔB�R���ݖׯ��R�F��
�&���I��ے��������"�������}����Avp9O�(��,i�  ��IDATG�s�ie��a�P_5�f��!�\O�:P�w��R(�-԰�!9�=����˛�wp���H���~X�LۜVy�1F��Y����l���dH7�S|�+�R�����B��:�D^9f9`�υ� i�L�U��6z��\oUڑ�i��ʛoLN5>�����=���iO
=;'�C�H��8=�x�8��&F����)A&@�I�Q�;@�rVa�"�/skv3O���d_L�HYخ���9��2�q���6�7yQ�%ߜ��,�[ڢ�� ůk9R
���axH���i�<��H�G�,m_�������D0��A+�XT�`��KA���#��Vts�"�2F�v�9� l����e�l�����a�n��k/R�i�D���ʂt�a:b�-�+j���I"���'E�(�	��cݕZ���f��8F��Y�;�
��@&]|��Jpz�+	���p���'�w�<K/�q2를8^2�����N�����Be�'���}�*S=����_�Q�ʫ(G1�GYG9׽l�(߀\��u��큺D�S ��*o>bw{�(������������bz�|5={����S?k�~w��һ�;駟?���+��^J���%�E��#i;rqu*�Plo��X
�P[��}�<�e����c-��ֵ*Tn|� e���N�T�il�?=\�K��������f�W=ɸ.��ի�����/�ڧ-����r|���K���3��/C�^Ca����a�ʩpf����R�2̴��}_,I'�F����S��rEC��=H���p9O�k@v��DXA�Ka�bVu5ҏ�r����;`�M��~�.�j�X��ۘ��;�;v��V��N�������	~r�����%�B�JHа�F�'�/�:����Fv9;�'_�?�;��*oNz$kF��"��������xZ�Ns�ci|t�J���E���K�������Un��Ȉ�*��(�|Ȣ��`�����0�)��K�N��F�� q 3�{�Vn�,��ŞL�[xw�~��.��V��P���495�FG��%�������ݣt�1dog��CR|95�Hrh�7:2�{Vn�p�w�NA��X�VIi�(�l�}��fdˮ�/뚝 @俴�$����O#�Cilt���1>F����/ۤ��]���3O�קqS}�Ϋ�#^�����F}3�ĽHː��4�^�g��ޒ�t{��7��؏�*^޾2���p�Q�6
�r�tr$ͅ���e&�iZ���}:?��Q�`�:1���k)�YTt�ʜ/ѪdRw��N�^�[�.�[ҢL��򯕎��,&qL >%ou��L�I��S�|)�2K!7х���W����b���vAD�2���-�_ ^
z�^�����v��lȬ5��R�h��Q��+k2��长�\^�K+��ir|���//���1'Ӝ���]=��I�c7]|A�pj��r�_�-T��QY���״�%�H����&r˰[IC��/k���zҴ��奩��8-�4�%�h���w��<�o�7����w�<k{��p8����{�94���}�� �l������B[��Z�!Gp��K�!�tV�LLYK��)��Ǔ��'���(=y���؎��eO���ě�G�ݻM����G��^�R>�p.��Z����3��kǻ�Z�NОV[�m�5P�����ka�@ܺb��L��u8	��L�g��D��܂\�W.�%���t�*������_'���o!A�?;�?ۋ��a
�
�X�V"������R|Kp�G�9�@@�ah�/�K�Ls���Hz�8��<�U�\J/�,�G��܄w5A6�A+g��L�F]�����@S�+��@8��*w������4Y��@��Q��H�o@J�"JFni|����>ml�������<9>���=d���{{4.j<ay 5_�?��ߤ�6 ��d��-8��,C-�ty퓽M��y��G���ڶ���У����459"<��>^I+��*�G��.U�J�9��D^���[�7�r�{@U���\�������&o%eg,�X&�B)�e�n�bV���:Jj#��~L8����owkB�_uP�[��A\�U��_���U�����&�-: Ќ�ɷ�*�V�6�b�\�-����/�BGǌ[�H�@���/6/�9��N�S���D��f�B[�Veq���>�W����)t U2@��UC&�D8�D�`�}ը�_����s~�y�Ν�{�N� ���ތ���V�Pl�����Ŵ�4��G���E��{�>|���'�W�l��#ͬ�3��jZ����@�#��➰w����B��e/e�x�x8�RI�_1|��!d'���kpLR�gҷ�>O����Rp����4:�j�*G(_��>�Mo8B��V:<8M��P���aό��1��[X��:��0{�Z3�f>w@K�n�!Ln���-�}qk��>��B�a��/��^���6[wĳ�j5���P���������>�jwk;�n�s�>U$Q��L�Wg�7_=L��s�O��������Zf��2�d1���Q�=˯��z-ل�˥xۆ�`M��3jB��3b"�O�2��2TL	pzF3#rɓp �圧������{�~]��w,�Y��@���������٣��`)ML��)|'G�J��oY��oy��4^�r��ɡ&t<
;�m��\ �W��w��=�Q!����ik{O�t'�h�9�r��X����:�%)�<�0�r鵾�o�yե*k�Q6�4YA�2�ݝ��P<3V�M��C�/��{`��<�R�K�*�ΐK�Jc�G�����l WA#_C�}�^ꏺ�����*u���s�da�Qi	�!O��S�l�3�I��4�}�e�PC��6=.�/I�*���d����:1U��c�|�;>>b��}ۦ�&Ҁ�[�\�ʗik�0moz;by3j����1[�L�c��vlBE\���Wv���q�Mѐ�ME(�� �/2��aƙ��{��´�܅4���5qP�~�P�����Zz��SZ_�J�Y�r����֯Fj0�?Z5�0j���Hgo���-�;a@�@��<wF4fx8R�P�u��.��xz�d�G3���Ϥ�ё<c{��dk�>���)޽�H[[�tn�0�`%޼���J�_nh(����k����~����ƿJ��|� �h�_��r�?u@��I���f��6���^a7����VS���j[���^�&���E::<���>}ZO�(B��Rp8��/�Ό�Gg�w�>�����Ջiyy6�)��s�1�>�e��-颏X��m%?B�2�j�Tf�/L�*̆��.�������.�����"m���C�Ok;ig��7 �Q�����l6=}�,������9�����̧Ry12��f���r/�k�lgL3R�YFJ�eL����e�^�}m��UP�m�-���K�S�v��$&&Pp�!2�F�)|,g�?��P7���!�����N�M��'{��P�i�P۠�Cp�r�_��N�F���f�ț��" ?���vhs�{����Τ8�7(�!2i�	4��O�A��bp�2��(%":D�-v �2]�"� x����<-�<�s�xM �)��9*���ܒN��AC�K:��')ց�-󙣋[���٤f�u@uD��*���� |ˌ-&�F.��poZ��Hϟ=H��7ieeQ
 �mO:9�I���嫵���Gz"E��`b+,�E�������3=2"|v�?�Tx�a	�� v�Y��`�v�5I`�㴨���e��K0��͎�o�y�������Z`�����!#G�W|���?�M?_���vw��t�_�2�v󍆚�%{��
m��BL`�)�p梮j,
.<6�#�(	�|�`q��k{zXϵ��@�q�fgGӋ���~�<�N��r��V���������Q�᧍�Oz�~��m��~=쟨�ET:ԭ���WH�S�Q���̏�����aȖ�\�����=ed{��`;���b���n���͠}�1������.��.�/@���N(q� �G�w��%l�����u��;y;�[�Ļʵ�P+{��>��N�Ϫ�	����IU
r�����m��/��A���FG�ؓ��(�g����m��9IP�^)��Ʒ5�!7����e��G鿾/��ώ��t"��q����PيҌ�w�g��1OS��idd�<sh���K1<==O{���a��C�Ř�r�<�>i��ɳ8���l�{X��q�+�E�RF%&��k�7 ߐ�m��gǞq^���c�z�e	!7ų*���8�z�.mox�Y�u��sχ��)�E����֤P��[���TA�W̪ה���:���c::��X�������Ó��o
BG�I�牠�e�ۘ$ɘ��Y�Rd&������r�,����ȗ-C*�-%�J�h�W v�@�e1f��Q��c�i~v
���
喧HB�hD���$7���@�%�H/���O��MTV�=1�Utp^	ٞ�N�4�C����u�x�6Q�.�4���z����x"��;K�?�~|����tv!��'�V<G=�/.�P������(d��(q3���[�Lf���!���8�+���ԯ'�ё��`u.��_���z,E~!�����z��b}�0�~���u9}ms�C*�$�4�p
�Z��u�\0�Bg`L� L���,a
�n�/�"��n�E�Q����v��i��LT�(��|�,=z����'\W|vrv��6���?�K��^��!}���������x��9vw0-*L�=��7���@�
�Ϙ�#��=�����ٞ�7�k��+���Ch�ٞ~�B��4�6t�d�R�hķ�=@��7&W�T�lv�G_���[�^�@١	9��1��X��Tʶܗ@)31�rk;�_^P;чR��[O���o]n���!+��2�t?��u?�r�1��2^�_H�F>N���|]FFs�rw�(�׊r4�S$�6�9V3%L;4�"�� _�)衤�l����S��?u�?>6����%E������u�vv���陜x��cxŏܡ��������h��mA��K;:�[ 7�G��e{����'i@
ܬ����Q+>�keJ���SGG'���u)�GzhQ}J�Ct�i�GJ]S�ͷ���tr��k
�5�ɞ!t��9�c�֠�:���H��o�VmL�4D[C�%(i�(�#9�.[0C�ߐӺS�=���f�*���ڬ_e��U��ki���/�l
	�;m]q�Φr�_����E�ua�	fLn��o\���;-4����Kơ��9��!Y͇n�3���tEc�iO|@���+ѭJ깔�Y��M�}�T��o� �E^]3�ɬ��?�������������*���-l��h����x�����i"�c+w:��xT~�'�DVT~l�-��;4ܓ��&������ͷ���iR�-ux�'��]N!��Y۟z����Δn�@��f�Z5fA[>�Ne�6���a.[� u';�*<��G���]��^����4:ړ>Z�!������c��%&��b��u�^��N��J?��֯��<��+>���'_7+'h&k���Vo���I�~?JH�U_넟�Hhe�W�!{��
b*K+�l:~��������T�w��M(���@T��������p���y;�]q�����s;T9=�K�.q略"+,��M�2�0Z_%�,���|0#�kh��;?;Ig'|�y)�v(��|���9��-�ܘ�e����#��)��Fg���[,r=�K�?�I��,'�<���i:��|�.�n�����rd<T��ƺ<Pn��9�P�����/�#�s����QO��Iiw� ��X^�	E��2)�d��El�3��f�C��jW� ���h�%�G���?�[x-{墴�����&�20��X��)�L�Oū�n�����>Ƞ��ce�{�$p�FpXڱ�� W�-B2��bԟH�]кm�e�Sa��XOY^��[�'pz�������`��9 � ]��g�(�v�*�$e̖�4�ȇHC��N�O��A%e�ڐ�"O�A�����4�������gj����L���r�\&�"~A0hVj+�T�ɛ��8~��R
ˉ�gI�4(.��z�iQ(FE��k\
��.����Mu�v�� �4�X�fI�3ߪ�B0E�欭�B�!z
ΔF^��2�I1�������Jϟ=Ls���5@�lo��_~J?J�����isk_�-����)�:�=����o3P.�TiFl,!�GY��Kx���U��'��~�ؙ�~����c+����b����k+���ϯ�߿K��m�	�T��a���%̜�?R�Uov)��oڰ��u�	<X�3x)q
b�K�ұ��� {)�V��T�^������<��_�|�\
��4�0���YXNա>O���[���ߧ?��e��>V./DP��kP*�Cq�<�g��U�[�8���@�v�jW
-#m'��D�Q��f��N��^n���ݢ���0��� �����/buJ�	�u�.hC��C��W��.�����+<3C�1n#�������VC���1��-2��1t��_�*f�XFt�~4��IE!��S��+Sa�>dq}d��#������Q8L+Y��З��s5&�Ơ!�Ԧ��۳�m�tr��4�t���S����_H�!�(F$��e�,��E�0�����M::��wr��M�)�0Qn���-����2�y������M毂b�E�;���AxLИ�|˒��Q)?l50@�d������C�z�q�H
���S�փJ���a@��w��vW�lC�6��j�+7�̆Lڂ�"H;T�^����2��QY��nƷ��9	#F�����J�:W��r�];�老�U:�Fz,�
]M�
�{�7��W�3�J�^�sRn�����x�d�����3s%E~
�c�%�L��i�`���<J�Dᴢ�p������r��黰EH)hҕ�AO(����L[E�-��Q��~��4>Hr,��ha�Jp�.<D�����O|�`Y��rk�Q�A����9W�^����4;;��=]M���R��-x�%D����~N���gm����{���ZA�	�l�Akq�^f%i�܍�1i��N��4���/]��`�1^�PDt.��T.�"\���T��BOY��}����Iz�0�ҥ�y���w�^K��o����ӏ��}	�G�3��Hq�ۓH�7��4�d6x.~�����s�@����W�&"��m����==g�d�0�ÇsRj��?���Ջ�>Fxll�B���������n����G)�?Ky_�R��%.A=08��|1;���$ ���n�X?r�\>�W;X)iG�݆�`�w%��G�	��V n���X��.ВwA�l�
ׂ�S�w��`ٿ[ ��ن����Ѕ���9L7t �+�)��pM���
�_������f�*9ٽSr��X^�ޮ��i8��b/H����J������$����<���d���#C.��ǖ��R~��NL����ae�~�<y�βB���T)������mE�da� ���5!d�k����B��ϺX���c�g0Sl�[N�93.ͷ ��]�q~�ޮ}i~n.�����1�(�����F�;���ȯ�7�˛>϶��!�X�ې3�T��V�trb�eIĽ\F���:Z|XL�8͌r������|�͉s��y�Z�]������N��?LgR���b`0���W�rڅLeN�f�·k0��� f���/�#r���Պ$�x����1 �������]&#ݬ���m��/�ʞS��s[�.&�oӥ4�NZL�q�px��ϕ:�C��a�0I��N��x;�({/���r;�����@��i���P�� "�Ds�
�=���cp~">߆o��NjkWhƬm5yaDe[�c�d��y����t�+S���CT���_H�� n4��x������2���y���V�N�㼒��ڮ��K����a3}��b{�'lf���eU�A;`�3��p&3�G#��:a,��0�G�W���͝S^~"*����w�榧F}�9��I��� �:��u(>wӧ�;iks?��@�f<��D�
(G�Q������!\�#�	��]*p炼FyY�?�R�onb�vbb�3�_�x����Ez��qZYZ�>��L����z8��,�O?�K��}�b{y���D�W�+� �m��h�o�3��p��Sʨ�;a���H�¼ޱ����*��fZ@I���K��\������A{"����dZEx]�u��e�E{l���µ��R�<�I#rI�nj:��0�F�,�[���:���P�,dQ�Ol�φ���!��\�Gg���ۏ�X����x�m���P_��IVfԿWVf��Ԉ?h�{vLA��{�[PJ�t�ƃ�2��~wx1~!(J(��q�Y�����/� ��9��Y�>�|�ppx���#C�7>=�=�KO�.z��+lq'�]*M�������J���*P7��&���H>�W`1�W8/)�]�����ړvv�k���N�	m �/Li�5�SS��������G3[����$?C3�����J���a�[	��}������j��!�R9�l���%�该>3ڭ�/K����9^Ml@ۭ�J3���5����(��RU�gƂ�p�͠��M]�|�.y�05D�Im(��+��?����O�l����-K8��5���	:��B@�ܲ_��I��
%��(�Ҁ�uU��@Uvv��
p��YTuCS|5LK�[��-�)A.���� �Ka!�����>	�1�R���udxP�NO��')��fno���hг���,�gl%����Wv2}U�� ��q����2�M���'с�y���YLi~~�������ٓ�8���zb�������~�~��u���/���gl�W��cV�������A�'_Q*>)�B<�ȵpX�tt(�\���fY�����e��r%m4���m$؂�LCFr5�/�s���[�
(�M�̖�c����@�7i����~�]�S�������&���d���9L'0���N\(�NX��n�
=��2�~V� �:W���1��xp�P�__��O;ܖl}��S����}�ӟJ�[�^z@c�;:ܓfgGҳ����������Q�,K�N�|��,04�
_tPv�a�C?�q��,_
� @7������(�W�=���"m�����5�;|��u�A�-,�����������/f<�f�������	1l�(��qk�#nBf��wB���,�Mp{�E?�wf�9Q�1V	[��5a����=�hăf͙���O�+�iqI�z|�3�(�,o>d�ad��#��m�[��y�o9�������MZwP:��+�\&\���]��v@q��	G��?ʶ���i+3�����s��\8:�ouڥ�KΝj���f����@FKl�<�ß:��Nȇ�zZ��V'��b��S�HD��8����aO�=�b�(I/`9�:j%��.��ڕ{ ��DiX��O�.�\F/`�Z��I#��NNJ<
<9Ǉdl�~%P��䘅���Rl��B�� �x}�~#}���CȽ�(}��~Mg.C��4)&*h����i �B���oA	A��gJ3�B2Ks..���M��d�����ɪ�U��N���A�M�f���m��n3��ӛ��������Y���vn� �J�׏]�0f�l��&��:��eW�Q��i�B���`o���:��e� ��,�n�ܳ[N�����rn�P�YU����ᎌ���2��0˱6,�F9U�2�%���CɒM�`Qh�Tl���5��R/f�~��]�^}�ͻ5)�{��%�Տ����K������׏��g�iN�����s�s>N�/J��)}��a�>}��lA�Y�2�V���V���U
�E����l����+���'DJ��DZ\�7H��F����VEɷ ye�6?�d[��mq��m�_;�[�6���?�ì��I�S���a��޳"O_\P=i���hZY^.��_o���.9�3���9f�6�[���oͬ�Ⱦ=X�{�=`�Wݮ���_eKȘ�a����e�˳aoq/�l[I�F �
{��: 7�A�@�Q4�R"����H�$Y
�Y����B:��R�U<\� w(�~"LF�-r��ꂑ%	|��0�y?io�u	�ݝC/�'!�-^�+p�]�)��ذ���[����!�'.Ғk@3 �Q~1K@�X�,���u<��a���l��������x�B�P'B[�'��������v:?e�`�����&;+��4�s�%� Y�"^;��k�.(���g���ê\�����C�vd�;7ޤs)�W��'O��>}����r�� ��4[�0[��[~�Kk�6�ؚ�A)�@�2�!���������##��(��� ��{I!�����&�m���'��|k���/�#�	T�s;yU���`]���@�xo�\���L��Jr�Mh-�B>41{� ������|�o)p�7#�P�������Dl5䴳(�m��(�[H��q*�� ,Ex�~����?�I?�����O��z��1r��PG��>L�}�4=|�,p\�|��N����S�$�U
ay0�6#��/�-�귃̿�1��R>�Tv}�D
��ڦd҆�O4��v1�>�����:|�13��t)��ڲ�o�\칎���ڛ'r������˘rp��P�Ԫ���[�X��f�A�1������,9y��%
ɇ )_�6�1^�r���J���I##CJ����Ә���H+⪲t������{+�x�����}���_ک�2�B��\&N`�/�R'T��w�B��_��MUy��~1��(�.�Bl��ڪ@��e@��a�f�K�wgjj[�靁|Ph��YQlY�O��b4��9���kl*���x��������¹7��:�F�0�m�iK����[`O�7�L>�_A�[�+n\ 4Y�e�V�{q��<������G��U�Eestɏtpx�޽�L�4�xI�����@f��{�5`�l�f�@C'*b۠�c"$�`kd ����B��r!۸�3�0�VV���|���c*���X��#����Cq�Ѓ
_\�A�glU1�yR���p��+Px�`�P<����{`;4��RV�nv�-��!�n���4���mP�ʙք�A�uAU�Ao)'�p��h+~wicX�e��hK��k��/��!�n!~9\��goh�U
u�l��7��L�Ͳ�c�.E��1�h��
١�&����t|����~��Sz�a;m������f���`ZY��[.��šA>�:OWg�꒏Ԙ���p�k��*�!{Ms��Ag���~(�R&-�
�s�E�\���8�{�K��7v� ��6��R4�M���Tz�:���g�⚭�.�p/��C�i
�/�3b�}���tkP�c��0ӈY3���P ����@�3�����1ӟ�O�����qS�n:9��x`p�_J������Lc�l�x%��T�����v(�a��kt���
8ReTp���%TH��h[F���m��B�z�d-r(0ڿ1_�P����_؈Cq�*��
�s����W�s�4!��[肴,|�x7���6��X���X�6�.Py���p��Ei��nQ�X��z�b˶$��R;7;�-hP��Y2@�&]�\p^a���؂�T��&	������y ]��2j����զґ0C�e�����OOM�ГG�������K��K/~��M���/����)�{�\�e��[>$hU�2�/d�]|)f��� �P`���O�}iQp5�����n~~���NLrHCb� ^��5�ۣ���VZ���N��rs�� ��bK�����M	y<S�
�tɽ��)~���$i�����@�97a�Opd72�b��>bQ�Q���c�]E��2ʩd���)|ɷ� �u�����s�Nn�!��Ee�l��F{�LD��)6�E2Q���ި4"�FB�"ˉ.���p�O��v�,�
m�`ŖPE���!'4e׳�Ȕ����xa/�q�ݾ����~~����z������1�9>ާ~?b���49)�-w���`��~�#�7�Ą��/�.;g7d�T~*�2�m�lȃ5���+�`b��Q��isk'�{�Q���;�S�Ȏ���}R�F��d�츿	�׃���ߞ��=<0~}�.Rz��� 3���P@�Hy.
o���7(R-$_D+#����3�K��U��0��1.Ę��+{����]��ַ�/������4;7,�v<��1&]�e	1L�L�8O�6��&�4t�a��@a���$T��io�9�*93�ݨ�|�
1��V��t��s
��D}S� ckܓD؛��n���#��vA�,��*W�piŸn��h���1r����|A�3Q��QA�&ʴu� N6�#����5�3�547�4G��T��KDI���.|��
_y��+*6��OK��ia����V�)C��w���T���ֶ��޾Ֆ�!�cU��8��"������)�����!*!��X�[�D�+xw�v�BEE��-o�q܄��P�,��I֣H��>����7o>����>��=�Y��M�$�I(A�'�lּe,n�<g(��d`��Ia&�h��101@I�i��I��3����pvfZu�Ƞ�]j�<J?��)k���z���Gf����S[q{�˒��`l�����&0x�
�rN���f���U�	8@ S:��\'�[Y�l���id��	��� �Q%ڎſ��q�id� ��s�ntwx���/�}h��0 h(�Md6����

��?���l����,I�6^�3fO��YU���g�%�%|���q�h��#cKx���f M���5t��g����[�������ǉ��ӟ����Û��r�(���Ā-�z�в�~ƧJ./M���Pp��)}dE�'��JJ 
"��y��Yɥ���6(�I���� �ҟ]�gyS�?���}z�>O[[{�������v��c�^8��7��J�aM�d�TR������Y�:/�m�a.S���1�z��	Έ�%p���\EVS'�����·���gi��C{�b˒���˴�{���mhs�@��Tc{���������<�*���QI�6sn����V|�(AW�^�G��O��0��%Zc�4n�V ڍ$��D��f�Uqw<2r_��?��{��L�]KXa����=��-��@��Zz�	�:���������?� ��^B�*�48��B#���^���3i�[���[4�V�EC����8�'7=�QX����4ܒ�S���_���(��[PP�!�P�	�b Vp�+��^�������]D@�K�$���	*��ˉ�_�Z���F���Z�����Ne?�`�I��LO/���=�ڮĖX*�;<�&����O��s����ΨgE=����ʚ�^!��f
�3�u`S`V��Vڦ��&�@6���G����<so��{��V�_�_/fϥ����wuy!���K_�x��B	�O��7����6���у���8����-l	�(���2n�חU�`���^�!��Z8��U�|!�n�jo4�Pn��y��d������C���dd��X^���,���F������wo�ҁ��H]�����ܰ�H�7�+n���R��AaH��tG��F.#��sX���C�\�. �l�S� �[[hg ��(�|9<���3x������߼�Д!�g��p�R�W����`5bd�P�/f��P\��v�9��VX2�
�/����/�n��37�mb@��e���*�b�X�����7�e��W;@n��S+*��c发��M�cV�qDg�:�'}[<y ������c�-ʩ�!������Pxվ���/]H�;=9���A:=S���RcCiH28(�у.!]���c�zz�zMN�dL�/�*���ܦ�B�C߇SO�؀J {AA�������GyD��Pb�{-�&�'�6mh�7�a!���~-��>}ZK�������/���{��Ӯ�@�������,�B�> /�E.�R^f�e���w�l��"�Z�0_�a�L�d���>�F��ڱN���]zvw�T���Pu9��ߔ��o�"�]��5�Nu�9��L�oJy��V�0�t�1 K� ���C�v�K���v�pT��>��(;��]�����R����(�MȬ
h
,��g�3�&m���^J���2Q9������З�Y	I��!�7���cuj@�BS0��q��-���o�",�@d!(�`R��!�	�r"�����#hA�N�A�)�7�3�Y���8%L��m�ύ�ܻ�h��@׻(�=cN�NUfnoX�/E�-����W�3R�X�u��rqq#%��[�|��vuַ�{i�W�� �ꯔMe���&�1�>�(5	@<�WA�i�^����+�ʒ�Օe�7�K��/��O;Vj779)��P�0Ć�t�d�u�NaE6�恰u��1���|�<s�>��N��#5��5�'�/�So���Ѓ�j�����./���
}~����Ez�q/��z=��������<�S'Հ�r� �@!	���	%�|9`(��/Ќ^�06�~Sڲ?v���*�<`��
n�S5dyд��7*���q*��7�,k�ػ�A�u�.��*iTi�B-c��'Gv�AEB���bǬ���-��e�K�(n28˖� �mA��_��naC����)M\��V_�uo��ᅸ;(�6�%��l	W��!�굡�uI�+!4�����Cv���nl��{��o����is[rJJ/'ZHOM{}곧+��㕴8�3�8�Cf9M;�Q����+�"�\Oru���K��܁b��M�'�ʲ6��>�L���A��q;�+�"�䓼������/.̦�	)r��.0%O���Å�W�vF{��T�3߹���	K8��3���<�pK�i0���ϯ����?�����j���=������+����_5.2����Y�b:`��
����v��1V�O�d�b�l��|�V�/�}��˭�S�A��WŴ�1��*m�sr��2o����[G �'T�`3|�G2C��p)����
�-n�C������2e�͈�҉�ni�Q���8s�!'Z�ю�΅R`��!8�y=������Z[=|��f����>ydx�O��<����n��΅�"����)=f�yz	rH���d��I���=����Q?��:�}��r���2�Q�:7>4@�#���l4=z�*E�Q�������er��R����~:;%=f>�l-tF>\��o8�Y��w@&��̣ӂ
����K�rBXou-�Ɠe�w1`���tz| ���[�=X��b�8={��f'G�Ѐ�)���7��:�뮧W�?I��_/rPi+�^���+�b��lڻ<$h�(:K7�-��V�2� O�]���s�4�6$�5��@ٸ=�Fu w��&4�œz1bW]U��(*��kG�q����������C�_e���o�O����N��tB��@] �����C1oH�1��C>3l�(�=��?:f�\$���/��AB�Nℨ�z�%7hw��h�œ\�����KO6��r���VڒB������A?�,XN�|-���?0eoﳓc+��688�@���\Ife�ֲKLE�T�@��Mܛ����}���2D�o��.>���?o;��O�çM܋;��XK̎>��0�����J�*7�&\� *�D���W�/���c����´P*��N _%��O�WɏK�Y�p�������{xx���[;���Lr������N�����45;�
����8]�AR
�+`M['����~����v�XC��J`a[{� ���� ��a��-�K�NPҸ�_��X��ۄ	v�ϱ|O�P?C���4�υ&�K�ib��3�Y�2#r�F���]�>�{�
w;���
@�Ny����/=���?!VE��FF��>�|��+R��g�<�ɗ��[��Z��X�I��3�)tbV�J���ɨ��٨�ԟ{	p͟��G�^�*č�[S���уU+�3�ih(���Oۭ�c�p���
&�N�%*���R@R��tn#-�Yu��� �r��y%(�a���z�=�Kie��D)Wi~nB�,Ja_�z��QΡ�%�����h�M�^}J��m�����6<�H#�t2 �"0�Z��sԱЍ@I�[�~TA�^ �C�u�eƽD���4s���c��P�V�^n�f��f��Qr^&��b�ĥ��GY�z,f��.����ڝ��J�f����ɖ���!X
�*��hB�;df�L�%�S��/�5��
%�f\�(���q�̡O`Gd���?�_\��o�Ǯ'�fv���@wJc�+�3��ӥ���rZ^�K�cCY~H��]s� K*��My(��[�hVsY���A3Z"���Fe`%R�ˉ�[[�N����}�����@cy;%��Ç�i���_��顃	8�D㛛��Vd�/�>�,�o�Q��!۠x��m��-�f�6f�)x�v9����8mlmk�ٱr+X/����f���\�dk7�ų�)�,�#�V�I��
H����&��{�p���:���V���
�C'w�!�/J8C��.�l���u�r��K2�%-5_��hbBڄ_]�C6s� k��N"��΄r�n���j#wbwm�z	�|33�z*��l�ι��$T6�����Pn�Nyr�/z����Ycz�k�LX��V�/�[���Vٛ(7c�ۮ
�GV}��pY��@�r;<4�%�ܮ�.��q>�`��M:O[[�Rl����s.���wq�6D�����B9K�b�\ ���-:��})��u"Q�6X�l�-wq,�s�Fı�O/����4;���A�Е��M��˟?�W/?�unhh����z)gȗYn�}@Ӟ� �3b��B�+}�B #[� *� /�<�"�B��J.�G���/B����_n������B��3-���������e��˂2��@�_�JAJ- _���{�J �h]�
�l�����Y�_��P)���$A��{����W�B�jΕf/4J��X1� +@Կz�^������~���nHfm��ݳtz�!7i`�7M���S���H���ilbDYݤ�s�ɷJG�R�1+�ѡs�.��[1U��E�-�3��9^ًG�M���F<�K�ݷb���Ǵ�����@ό3;'�4>9,�v1=��;�qkhXJ���o��+�,�*;㺜�nd�f��J�Agŭ���tK�*(��oy�;��R>�p!~����go�LNV�ɞ�KK����)�s��ڇr�ēr�j���,�B��7�l�mA�i����J��u�3V���.W�gĿ*!c�5�I��\SA��*{֍�r;ڿ.}�X�!��#s�-��S����Ѐglg�&e�{��<E��^J����%+�x����q��ʂ>�FX�M喡xaX��o;@���D��A�.r769�pff��dMOOH�e-������֑��=����5��b�my���Y�
6�\�ݡ�-@&B������0�%��1S��jחg�_���D���%�L�yI	�3�(wv��Ǐ����u���\�KG���A鱟����W��0m ����A�[eV�M����C��2+�+T
#��h[VlK��=X���oi�� "��P��+�Uy�+��Rf����+��a �nxo���B��G}b�v��Kd� �YQL��=W��B<x���vhhR;�ϡ�1�fAB@#� �V�ȃ�`�.��O�<�w��~�����gR\y�6<«�Ѵ�:�K�E�]X��Uh�2vK cI:�)㊰X����fL��L�u��`ƥ�*���E���M>mH�]��{|�:PXd��蠏L_��[�8��;��i��rr�e�.r��o����*�r�PAT!��M��*�"gw�q�mXd�&�&���s><L�{����q���K�3�>;;�VV�#�����Q�._A*�s��1��
q��
�i���o�e���*.j�4>��
r�wE�Jp:���>L�LVn��&����ݝDh�F��@Y���Y�[`�:	k9�(��	VSRn���j�V}��Y�+�`�8�2�'����=���s�"$?�VڊR��uU�3CU���e�v�tɤ���	�X��%�,���Q��L��MyƖY]�({��籞�ٿ�����ŵ�aHe8+��PBӯ�Tfl���nP�������Yc���!�<(K�B�f�Y��GdCr[��N,��WҒ���a ����~+��Ӈ��O�W/n̸��np�s��}r��!��zk`q+��M�(��4�@����CB�(���yeG��<L@*Bߩ�-D[�z����6�7�Q�؛os���r�T��3�K�&�{��}���$9�����9,��N��F�6I�C�`�ԓt~vdd��*D[-
.m�`���/U��VL���ڱ�(@<P�|e�ԡ�Q��ްG�|��޾�C�w��5�2N#�tYb��0�?YL_�8=}�*����-�,]�*�]Ӆ`�KQ�`�P�`^5ʷ\w�<�K�9)c=����4��s����������D������M��3��C��Y�t)��| 
.t��g)�B�y��)��;�6��!����ҟ��ThY�e�eA4�3�\�����ﭾ/�R��7���f?_fo�x�e%ԛ��(�X���{耶L��@�/<Uޅ�r!i�x�/h��P�4¹DK'�_)������Y�������$��Z	��6[nK�����%h�:�g��.�fzu�@�9hG(J&�[�	�dV�W�|������OCy��cm���[f���<k�t�g�:Bc�]�h�B�m6*(\�Sʤ��{�^��L�OH�e����
�/7�S���u��?���9xƾtRh�,�! ^�x�g��|:�v��k��,�]c`�Θua9�S����/[�&F�=ѣ�r������P�dXO{x�r��޼ZK�5�mm��X��3��VXS�S����\���.lB�����L��W0��	!o��O�i�v(����Bm�&���yoN���
�&�f���v�-t`�m�1�>�ᒡ�׮��MSm��e�e# U���7cg�]���#fhX(��݇���������as8N;�m����[�̧�������'�-%#Q�ҷ/�G�O��V;���GL��|d�v,�x���"Kx�"O�K�m@��!��50���.◰�]�)+M��>/���;I>l�~x-��׫� ���Yޡ�>}���?[M++s�
_��VCV�@�nC���[�٫M����2~��Ge�X��eo�������ݧ��{�N�/ӕ³�vll0�\=\L�K�����<1�y<"U[�I��1K�Z��A-�AO'l���0��/�吲��e`Pcm�g��w<��[7�>mpdd@cִ��NOǇe����jҒߞ�*�hCwa����\F���;�?�v����/�،@��Yʸ�wӭ8U43 %N����d�U^e�$|ĩM��D^}O�����D�ZrŻYaLOw�K�
���|�{�e���q�	a<�7 �(�4���b�i0t��߅=NQ�=�� ��95�@�AS���
r� |:����$�*�:��$㎙�r,I��?�-t�J�_�]�I)JO����z��!),�9<�I?�D�ׯ?�Tf:G�&����󾒠�@I���Mg�r/`�0�[�ۊM���Sp�g�T��y���:�׉7�g�OJӈ������7�ҳ'�qa:�JH��ak�"�}�����Cz�W�'J�?�s:�����b�gic�+@��[ǫ����R�j3�j38ޗ-֨Z_jSg��Ǫ���/�v6}��S����J���@�>�)������~��z�~��>f����� ��
/�Eچ��|��C�Q��vn���pi;PL\UH�c��Ą>�M�ae��/�����V7#�>]mQu�(�ff�5��Տ�v�ճ�3~�%}��9�\�Nם��f����{��T�.��O;dS����iY�p^BL���1�6һڒ�H�-�[I� }�/P`Y��_Px5o�٭	.3L�ghbp;"1�W.sE����P��wE:O
�FA�a<���J�A6Jf�ǖ���Ҭ_OH�������YbW�[���[,�(�;id��{f�a�M���m�9<ai�4r��˭|�O;dy���i���U��8��#����ͼI����}a9����T�g��<hSndR�+�ٴ]F@�Aʥ�}� ۑ+aF�d4�/�@�P r��}!ZO�{��꒷�D�e�3�7�L��������A����4:!������5^�$�i�v 2놊.A�>�E G�E��A�jVv�>�V�v��:3;�u�sz�b�6�U��E���f:������[Q%��ҹ�NC�� /Z_����E�D��6��R?�dp�8�Ѳ2�M�P@��Xʜ��W��򱌡�8���H�6a�3���K.3m�ߺ 4�
�`@�e�$�}�4h�q�=�T�%߈�8�U���d�����DeΌ��(g��S��?)�:�6Pn.#�r��
e
k�v���^��|r�Q���S���8��M�:�+ :�Y�+��M7��O�8>�*x7T?���k^qp��,��g��M�o�,G��=I�^k�p쎆p�#2�.P��$
G&��ԑ����� ��m��ǌq�����dE���'���X���=O��9+��WB���қ�[��xo�H�����5�K�3�b�PW�
8p���f�#�
�ut�1�Ja�|x�Xp����Bz�h5=XYJ�R %�Q�/ί���IZ_;Hkk���9:<�R�R1e�C�˴�Qg\�����2ǌ�v`��Y��j��"���`�G��W��7i||@V��#^�>J�������?K_}�(-IɈc(5����[�Ц<��)0����[�]�s�k��tî�ʇl�Xɱ
���Np��=P��ܖ{#�̊�6$����n�u� �fi$��/�{╼:^B�(W��li7���&W��\2+819�>ZN�|�,��/��Ӄ��Vx��jo�6��a��3��0�%O��\��^֠A=^m�n��L� �j��B+�Q�?BB���Yo�қ7k� �eH��J���<�>\�G��SR���^���Mc70�P��8w�7(�������e>p���dȽ���������C���HY3���8��	��ih�W�/Jn���L"�(_��5C�L�,�&�v�hb
������ ��
�N�R}�+^�􀲽�g<eK0�V0����`a~R<�k��b����v W�"j&�99���M pAڗL�7Dؚ����D��B�ʲ�;���P�l����d>Z��A���Rǭ����/�׃��W"�/����7rf�q�r+%	e�'���Q+��D��R)H����*|��!��'Aɡ���bX:Q�R��Qy����;읁�/��&��H�B��d�=���pR����j�ʆQ��/��,��ҏ?�N����@�������k�D��k���,,Jn�7�+ R:�C s.��9�,"���m��$���r�Gؠ]����~�Ԝ���>2�m�͍}z�@Ae24̾�q��2Rh�Y"fx��:	"�r�U�)5���%�����xlis"e�2ML�%6������i���N�wߤ�ﾑb�,=z����>�w9z�����72�6S}!M������Jye�d0��E����	� �u��
ąXP�hc��mf�ȅH�� I��[�}P�Es�]�NCa��ys���܌����?|����]�߄��W���GiuuA�r̯���7�N���ˌ�-3�V� ��g|�Ǭ�2�� �Cb�]����'���a�?��>���o�8:�����W���.��������Y�4��|)JK3izfD2�W��`v���	aQD���[KҤ[��h�!n��a��>���K/������ܮ�3oo^a�����|_�L��irZ����X�*1�Ο���8�-�"��+�r���.,6�v傫�'nM������^rd���[)�|���&/������`u1-ic�
����Ty���}E>8,��۝+�Lܭ����M����'�g,�:�������[:2O ����A+��
�v��n�e�
3����*���X�E����)���5������B�����q�(�E�-)�@V�����C�����D�Nh�o�y��(�qaa6�L�{��5���u:<������zz�~M�� ��]H��艚��Y)SJ��\b��MTʛ7>�Jܝt�I��c�Z�3�ԏ�(P�c�d9��56�ad8��	�у�$���Ǥ���hΣ��~�^�\K�_�i0�7�<�
D��,���>��4ʧ�؀t26˽F��2ap�i�KZ*G8.��H�=z/=c�iJO�.���z`|����sRj�Ҋ���6n�13�³�ڒ;��.�v�KG6 ���x�	����/_58���+�(,P���&WŹ�g{�P�"����v���a��8j>~]̖Y��a}�����Ջ�j����������d���ʒ%�M�g�xE�[٨D�$_�J��r�xFy�}��-���0���>ŷP����ٵOXdw���=?����@����0ϛ�I=PN���a�He-9�kU���WM2��&6��4Z���j��V��T/�����Oے��&�p��v���KR�yC�˝�ұ�A�$(���}k���w��	$�	Ey�`6�KW�3`���<~(��׻iccK�о��S�)�����A=�L�ò��ِ�&'�[#��t6&%��to�LrkdA������ ���E���
�ns_w]�RR,�eo<�����p��PJ��ʸJ���S�G/�H%��Q�8�a���iQ�$����g7�@���>~���ݬ3C�0�u�LCn��:w%w�ބ�08M��(���1;��Q���銙��)���3���?RA���������<=3 ��E*���-�wUnR"9��'�+S�7�� dEWa�Lqǵ��諄c��pd,�<�v�0�:���i��>\YJ�(}�Db:ؽL����L���mz��C��;��4u�:W��aX �zUxʫ��'����bo�(���Ci�ݸ�����Rw^.>ˬ��١�'���&Ӌ�+���=N���az!%waf8�������}�u�z��R[΅���ܗ2�H>�?L,�@ٻ����D�TuO��I��Pʻ�_�g��]pmd˧c�� Q� _#�v,�^�wa�G�(�:������G����j}R
cݣ���o�?�����/ңG+ifv*�h*}�<I ��M��&���'F�y�β��I���K�[�o��ѱ4:>�~0�v�X��޾ݐ�M�G�8B��4�'p$��N��)�SR��o�-7�Y�/>��u�C��@.��y�ľ?���Ѣ_K�J�L�㧍���'��Tʁ~vI/�~uρD��%MH�.���.��NT�oc�n��/��g�^�r�iAk�r�.�hc<B������>�˾�m�H��76<��g����Od��.�m���u⦣�3��	�+h�� 8��\.�p(՜�j��=�z���(>��ƽxz���k��ڀ*@��P�U�?a�y�_����
/x����P����)g^g�6Y�֖Y۱ё�ѼJ�|����$���x�D��1֡�t�OaB��Lg�DC�rz�q��9���z��bCygm'3�<��k�Xk���Q���N,���I��Q����B^A_���[�H@<8���OE_��諂�hD��a���Z*����/�<����K�3i�]��wwϤ�n���^���7�/������8��PnU> d�@�r
�:Z��,�L����-�Pp6#Y������k�uvfL�̧���gOW}�����?�����9=���Յ}�fgP^^��:[�@�����uxc�� ��eP�"�@��
�l;~�y}	��8�b!�� �)�1c4ʡ�1�����J>��^��N�=�L����p<�:&��x���M����ՋG����[��m��D�ΰ%�a�t4-��О�@�g�5��\��v��QbDq�CuX�p||�#�9܁	��~�������UߛK�Bv�`�j,O`1d�����(����烸RT�R/�v0�z���־�-���2���I�pػǬ�,x��x�ƌroiC&��5|.�%L�N�<�E��|��X~�BH!v�`��ⶶvbB霱�ɑ�qb8�24d�e*�{,��eS��|2Ma�K�����B�n� �&��J/��o�s薯��W�H�]|���ҟ�^�� %~oY{��(h�����N����K�ې	�4U�SN���t��f��UH�j�1K;�dD$J�P2���Խ¢uPج塣�ΰ��;��򂭱���nppK���_O���ip��|4���ƍ1 �m�����ө���+�ɴ i1�x)�#�^o������Eykm#��	K޾�(�"A�E���$4�Wo����*/f�=s��R�{ȳ,iP���?z&�ŗ�R��t�1��嘙`�ߓ�������42D�%+����ަ�������K�@�C��0�'A*��J������-evq���l~(�&0��O�1_��e~(w_t캳G<f[o<� ����6J7޿���\z�d�ʭ��a�9Qَm{��c�vtt�t�H��Lӵ�`N[�<� ΀@�P�!K�( �&�v�
��W֯�+�ؙ-�@Z�=[�h��*�~���v�����ϡn�˶p\)hɧ��C���>�Y���G�{�(L,��䨃�#)�>I�1
��aͳ���ų��ɣ?t2#��,��E���+�L�Rb�x�!�0fy�1�a�M�b�WU�Ж�Ծ�\(�1DST?�_��Y%%z�tX{���=o�������y��'���t�Χ��8���[f;�>Y��+�9K��mo�����7���K�Q�'�(>)��	=t��'��EJ�=gi��S�|4���Rz���Ƥ���| �)D�M���Hf���((�,�v���!��*;��h�Me�Y�Ӝ�Ʃ�����63��YY�Eư��--����v�b�֡x<�I�3^���dҍ�BI;���S�:fvo���5�4lLc�F�޽�%Lڒ���"�b�?j;1�³�̢,�sd��꒺'P5M^w�Jũ ���J��։! ���D��1@��'����J�8e�O��-��
�R� n�
����Dx����|�Z���������
�p3:а;p�^��cew�'u֢�ܲw��|�.�O
��7����	��!0)��n�,�5�UK	����]^����7��qy��L
T�_(M,I������3���b'���U1��z��@i>�e�����[yѠK�� N5c��� ʂ�<P��A�e�=�(#���R��V�/�ɱ����lz��Az*epnv2����]������է���7;�P>ה�[�٫�U�7,M��ڥA��sI��r[�!0�[�cW�q�2����b_��k)�inz\��|�J���'���\���,��@���%�����������Qv�`eJ���W�B�?U������%X�2fPȠ?�A/@����]G�� _v��y|��2]nC.��,o!�̐��+CdTHí�Ž�:��3}�0�ep�[םQjh�B�hy�(fIT��d_�D)Ѯ�`H�`Iχk���OՉ��7�
��'��z8[NO� .-�O�Z��%�������g����ʗ�Zh���\��[
��Sn*^�)E����^������fz�a#�o�c��O1r\-��/�&��b�_��%��ʭ����W$x:r��ڽ����ɯ���q;ʡ���z��{�v��+�����3����ZK�c^�AVbY�P�.����]^�o���&���>��@�ǀ@W�;y�.���tYf��r�q��	;�i[u����E�-oKQj''�c��a�B�G��]����^J���V�r]��-:p��B	�=�.�`V��~�n��+\��Ý�t�f���"�� �r�ɱ��k�'b�"H��$��'���m��bD�kK������Í��>lsiP�P2At�=�H��J�EP�.d�DO8lPo��Y(*�ƣ��
 eb�wD�pF��0{���`$n�͈��6�
O�W�ē"�T4���m;MӪ0u�@�ұ�R��B0:��q!\ȟtJ�0a�ʡ��ZH&�#�����ka��<�0�����_���L���/I��9N�q-}��{o+spx�<b����!�����@wng%�J�Q�W��TumP�W�K9�P(^���2��t�C�����.���`�����'�]a�4��������_Y�+.5to��r�}�� j�� �^B�2]@�z��\�T�\��	��6<��_D��3ye����8��H�N�|��_k?{�0MMN��p�<��_j�:I��S������n��;4����%�f:|�7�=�nx���4H� ��\�~dU%��+� ��̞��}���~����c!��ۧ����;o�4ʒ�EO:;�I�[W����������?�No����� ���8��,�L�*he_�P���� �U��Q�hs��f��r9�p���O���6��k�I�Fqh�����7"�V���_ i�6�-���Q���9���)x����6t�:B84�����AFe7�i��HBW��P�M�mɔT�0a�!��o@46\�)���L吼�޸&o�H��	���8�ٿ����ҥ��$@� u����d�c�G���2$��'��
�y�؇��(����t�)��iZ������8�9��.����d��q�����
��ʴ��r^� C�&�vA�!�WV7��?m���ܐ���K=��/K��G�<�97;�:u)RG�JgǧiG���-�g�k�� �y�R�D;k�f�P����,�-W�0�ٱ�	RV���Q*�"���i�GI�h��QU[�V>6:���y=H����/2=99O|�|px��v��O�uF�U��{���_���VL�+������#pk�0��J�(��CH�U�W��A�ڏu-�J����?�Q&!]�9J�����s�٬+�����;i��Z�o�vU�A��R�r��%7䣌LC���m�?L	0�
�6y��j�ߨ�Lf�}n�Ҥ�q�5M�`��+���?���pf!2ǉ����dWb�9\�w�Li��5djs�a��jȷ%f��_���h��Z�BP���+��QVe��^�K��O�R����9��{w?������l�O�11K��WќAt�
�iq�"0+9ݒ�kL�V�2�xK#C�]�r�����|T浲
���;'ic����RlyU��t�B�6��IX��_+�R�-�2��	�FXڱ"Ԋ,����	�k�x-w�����R�cieyN��f%�y��H�"���*m����Q��L��b�e��BR��P X�$��������u�o�M[iMQ6��\D���9}nɋӑ��K�ߜ�A�;51�V�f�W���_<N�,J L�r��-���ӻ��駟�ӏ?~�[���T�u�j��*O�P2�#�C����~`J(#�!2S�Y��3f%��o��v���/�7=Bz�&:�lPʟ��ʦߵ{���^�r�Q$�4>#J"��VC�<����ݛ���s�V�qe��P�d�+�|NӇ�����||��7��6���؃�����PZY�L/���M?�C�RZ��J�RFn�`wyz"��Y\�]юR�1���| �z�o�nnO� ������C�+���]pEK@���7'^}����X���w�N�JK}�C��wiy>��J��O��Q�a�~y*�`�c��UP��@"oA#�g��q�HTY����a��F|+�7!��a�[^PI�3��7��~a	�����0���?�ë��0˨�
�`54�$cy�G<��I7����1M©?��]���uvM8�Cǅ�/�p�'ML�������J��D��G%�����V� A�1���qu�D�I�]���~J8�t�}N������tsX�5�Vp��i�Z�F^ت?���WD�N�%n�n�-2}�;��)��.��E�vɸ7�r�(���D�hX
Oi���f�IE�M����7���)�8��K�`�٭@�*Q��	��iH��`ҭ��:Z�:�7F���ko	G"
-k���(�U�Q:��A22�6HS����E���|/�����O��/���=�y��?fg&��xr"�vji���>܀�`8�
�xz�R��-��ӎ�"L
�~�e���RP!���_��i�*wd B��MЍ���S<O���)6����lQn����H�{)�y!)�B+��U��V�p �:�z��P�3(�#�H;��$ �G^����!�Kϥ̤Ag�����yz��aU�x !ɓ�\G�ަ?����N
�0>��#��z�!�ӳ�)�~��,��a�G_��߿ (�n
l�M�?f�r�8���M�6��	H�>,�G���(��j4zWĭ��=��ʧ�s�@��p	(�qg���/�~���2��Q
�W��?�J?��^���8�Pʔ�&���8��o��o�M���W��l��&�K��V��#ugdo��(}�|=�+[��&G�CG�+`)�Htx�������ol�7o?����}�!�q�,�8$ N|�d%-��I�ӓ��&��u�|"+�U ~����㲇k��R��S>,�}^����Fz+���6ӹdz9�����Ӣ��i�52$�E�8���
��/(�xj`�n:Ź��!���f�4��7�4㶀j%Qt���B��d��Z����[��R.���=����9���.ں�-Q8sf�] �vo'�?���r@��i7�*���#ٖI+�6K?v�v�sh��cNuO�D��H �_�\Cu��am��T�d��X'�%�Pase�g���&���ĠFCUF`�x»St|<�?(��w�)"6�� ]��IN�f��6y+`�Fؚ|ȹ��J�A_$�rmp\����_���/_mr-���z��9=�)���DF�\��|H��	��/�H1�oԡ ��!��@)���:;�?�����Ԛ	��^�7�U��~���Aj�|��p�n�S��4��E١��c��|H/2� �A�[�\J����s���r��c49�qzZO�#�y��×��˴���ks�'��	�ʝ�@�+\E~�
2�m.߀�^!e�	#N�B��P&��C_/
���Uf۹a�����jz�p��}������O�{�z=�|�.�{�1��9���<y'��aOŦ�����2�4dz�]ib�;94��Z��+@���q��vo��.!A����ҷZ��ʘ�~�[�Tk��A���Vt����_{]���/������x��v���H/_}H?I�}�f]Jǡ״��+�Ѵ�:����i��g����Ȭ']HI<L�g,��O�AN���Rr���V;�,tؼr�
�>�=�{=k�y��7�?J9ԃ�JO���lrjDJ�?.[\�Q|�d����f�6dZ��Pg�m�n��n�Y.Bc��v���'~�����t�̢YA����g6��96y���9�ǌ��h�!��?y�9ڊQp��HM,�~�	Dr�6�6���X����;igw�cT9� �LƷy�O�Y�?�=����Q@;����S����B'���j���St|;��Q�%L�[��Qf*,a��q0H����E���[`����$����D��)d$�O((��I��)h��ɯt]�`�5��˕czpVڡl��>
(��d0��(�&�6Cv����h�=NSX���Q�xE������466���QNN/���+��kǤ��!�5�6LN��淁Uݖ43��@ hr�V����|(�&�sieE
�¼��	+漉c��])������txx�`h�z,��f���}��L?4��(�V4��֯�!.+�!�-|��l��_�d��Eη_J�ssl#�!d�a�����=��)mln��뫼�C�;Mz�L�g�������Z����:�@ώ��e'�ĩ���kl�t�x'�����2��>[M�����9^&���� �����O��]�ӟ_�7o>HY��W��z�����ʐ-�����������'�6���(�Ff~�/���e(�(?��G��ak�����ID�z�E�6zW@Wa'�o#���,iwu)��<2׿�3}ak�5D�A��f�6����$o
���n�^s���\@Vl��"|�ӕ�gW�~!C2��P>��L?�$W��ݶ��+���48ԫ�����	��>M��.��I)V�j����!K_/�P�<B�q�Q�_tt�L�m��1H��Y΁a��!%՗�����~z��mz�Ꝕ�#)ݴ{��>����~�\\�U\��!�[��ܭ�6h6�<;a������]rp1�/���f����ز��E�9>��_��gR�YvA��8���.jm@��V����*�&���M��OƜ�/��d(c��Pf١�5�GGGnQ�<�H�����&�؟~j�J/;%�Ï�K��W���*�&&���<.a��Q2����/΃gY��yv� &�#�m�W����˯Ro�tc���V6 bGB�Jm`�8z
��҉���{ �&*�.BC.t�%r��D8.i��.@�*����WѦ;5`'i�k+�ӓ^�966*eH�L��Y?���qOƧ�R*��(�������F�����՟�	:<J���3OԮ��B��`y-5�8������L��^���&�,� �Җ�K�m�>Y(V���unX	�g,��dq<ñw���S0�R�������)�J��Z�!��N����a]��H��,~[�!.PY3�m�F�W��[+�r'X��h��W�HR0��J�����tz����㥴����q^f)z���m����^��~�/�}R��d@¼�S���+�Oe�2S�[��Fe�j�]D���g̴���t��t�}G�n���p�����K;��`wC{�|o�ԟ
֤��~�䯀�~�~H9�-l�R����~�=�\�ȅЂ%���ʜ���h5��?=�N{z��P��o���/?�7�wۻ�锵AJfد���ʃ���ţ���Gi��|��;Ӹ�Xq��a����+�Z�6T~)��"���+�_2�G��y����^j��}!@�0N*[Z��r+�pb���zؾ�R��+�B�*���k�ʊ�������Y���Ύ7�S[fIo,]b\��uv�������ݴ?d+BO�05*���3�ԍ������s�6Aჿ�������m�����/�F�o�Cjkcin~�1�T�m
�����_�Q΢d� Rkb��逺�ui����BI�����wBM�i'�M��I�t�H�
(.���M����L�_�V��1J��-�JS��M�h	C8A�q�����FI�4����I1�?}����M�@���ff�C+frt ��:>9��`��(���N�r��P���8/�!fPv�ї�ׁ���{�b���)���ӱ�5�%�gig��	7�J���KTPUgi��Y)��$l�l��;+�W*�@��X���D����9`���/4X�i��K��K~5>1�Y̳�����>����_J/_��6G�G�e ��8\SA��F�����p5�F]���ȊmsƖ?���i��x�mi��~��4���{�{v�x��z�������?��U�o���Rn_�#��ӫ�'E~`d8�f��	.Pjɛ/dcg�5y���5C����k�}�{��<7���wr�ӗ �
:}�;�:a7h�|� X؉ ��_�,Z��J�;d�L��7�W���&;W�P�����Ѧ#.�y)��o�GdQ{���_�?l�?��:}�����#Jb�J��r�����ͷ�ҷ�{���x�ff9���]�?��ik�2��4�#��*�{���� ��7�8��֕��=���O����F:�;A��
 K)���_��J�2���K>�������۠3�eD�,n�� ^�K>}��m��J���XS|������=<�#8u@d�ݐ�`opv���J�-���E��@�Nܳ���K��Є+X�=n��M�X,�T�Ft�Y_̈�X|��,/!;��I�SQ_,M`+O�>�T$����@�J_k6�*���9T��ʧί�eG0��(����u@9�
>3{ #l�g��n��E�Cօ�M�c85�� ?�������fp⍢p��4�E��ܳ�a+{�1�m�ʮ�	���GZ9�P�.���W�(���g�W|�䏓D<�-gv�,�}���|Y	"i�D��
�%[�)����h�|�A��AH�'������4��Iuz��+''d����㴫�}[^��xQl(��
��., =��"�dr1����Ƅ6���`gF�Wf�{ON�x�siiN
a̰�II�р�qm?�y��>|XO�{�~�G��V0�X����^���]��R^+��S������S���&N@�>Ӏy�&5�,-N��OW�c�3dF8%N�q��KD>��(��㻴���\�Q���ŏ�"w��Rn��A���.h䪔�F=���r��f��6�$\e�%��xݠ��@1�e���ao�ВT�h�%�L�ȹ������ݗ�ڱ+=��;�l�+���g�zI��3s˫���a����봽s�޽�L�^L��n��=)X|�C⃟������b��'�o��Շ�ir��'��\p�d�e���+}�n���?��E�Y�~��>�}��zQn� �C.$O)��)��.N�D�T�c����{%����Y�r��:�7_RDQ�\���f�co�w�Q:R<K;(��wf��oX2r!��(mm�'��2bR�������Wl�����/�M(��薂Ľe�yi����٥Fl@�Y<d�cvW)�7C��ѩ��?8M�:Ǆ��߻ZLh����&���m�/*��m�=P
�(��7�i7�W��g�I�\f�-D.���!��a"AdY竂!�Rrl���I @���akΛ���U4f��e#���h!92&b��"��i����P��<��ƕ���Jg4������ ͘]�R��s����۷�ЛiΎ��^�c� �R�r�R��M����C �W��9�LB���gg���7%%JO�z�+Lf�%$�S�H	�e���_n�.Ӑy¡������>����S����R�k�D�_;K���6��9�2ȇd��p�t��c=����?H����rM��B�fZ��k,W�~9
eJ�yv�<�����Pęi��L�4�=���ɡ4??�����$m>��M���G����|��
�j%.��5��
T�(u('hs�\6Mh�/�lQl{�%���`ҟj�|���OU�u'�C�&�҉��ڧ]o���?��Vmq`De��I��UV�	��@����߲��x��5¨~N�"x*u	Oa������5#<}������3����.�;�����q?�l/4���1��7�U�X�a��2�R��$��@���~�_�MZ����P��̣��J������M��C������@��>i�,	�B���ݣ���V���������^�?Da�N�j[�#=>��ŋ���=O/�~�U>�:=�(\>2;��[1@f�,|)�����Gz�o7�7}r�S�Rn7ӻ��icS����o���c���'�RΗ�8��^� �-d�Ȕr��f�G����e�Q=l*C��e�� F�g�G}l��=�}:$J�y)���ku^�)Ƭ�������N��J�����9r������ӣC�"�{�1Lix�u��
r]t �1��_�Wj*#c'�"�:���!Y�ј��r\qR(�q��Ʀ�w��x��z��3�,�ol�HZ�/��E�5��C�i��89@�E�I��Q�^�q�E7��ί�NY&���+ܜ�P�>����L��r�u��a��\!����vv����Y��W��t�<��?��mI�<s� <ܰ�G!R�$������S�Mh�5�cq��v�t�WP��Q�V�/��L�1��a��a��p�����	Y������lC�����49ɒ�i�n�! _�i���_?������
�_������_
%�蔁j?��>�uN�����e/��}{�6��ıN�0N^����z�� A���s'"C�B����K*(�3��4�	��G\�����`�B�Z#�/xKH��*錓��ӺZNWC�=88��士8�,�t3VPẍ��)À�`w�5X�йuY�\J�^���{3(�=��g��3���3�������E��8H��؂��������\�u}�F�_xp��y��bk��!�9�CXs�鸁�	�a[�N��6t���ގ�>�����>h!/�ob#��[؈S���,�i�d �:����@��S1�_��+	���EzO�A�W�(Ql?��7�K=���l���~���>�~����mϴ1����ieyƊ��gӪ�3�/�v���Tʭd3����Rr��ՠ$b Fِ���[)��gWik����w�ioO�H�C�����hz�`I��f�#P��@�� ƒ(Ԡ1�����V�G�
lo�mC�;	�=�4 u���;v�_���m���v��ٕr�
����<I0;;.���wvrK$κ[+��?��]P6�t�U8l�g�b��b���r-x�7md���� t)�~��чj[�Nb#�YN8&�&&�<�3<<�4���ĉ��/��o�A_�z3���J�A��8�h/����:����U4�X��P� ��\\U��r>m�rTC���҈��*{&�r�?�L
v ��'�K��\>�k~v���r-��Hz���6�=�"}^�G��?�VY7�nVݯ��`H��Ѷ�����w�	h�UM,��(a��b������@L����$з�n��J�j �)r�9L�b[�<P ӈp�f!/�Y)�u�&a�h���(��	O�z@d�Lڠ.������Y��a'}/����k���8�2�eZ��|A��+�l����\-L��N>�i���+]�:b��R��@Z]�K/^<N�������c)�q��Y���v�^�����ϯӫ���1�+_�� ��j�m��*��lVhco�� QP��S���uv�Bp�5��b0�5�*e�8|�8�����+ⵅ]n�_2�ƨ_0�S��6�>�وSŻ��[�
r$�%.��}�ֲF6g�e����#Rэ|��Ǎ�������d����g�Ō&&ؖj�S>~Ĳ>��M��ܢ:���[�y���ڿS}��4xj�.�#�)����A�=�~���6����o�a�[i�F��dLr��b�]�܌g<���田K)���e(Δ��ՠ��J���@f��k��z\�t.e��Plwv��)ߊPg�CՔFF{�6��������p��l�����Hī����8�;˅��_c٨d:��.�\��T��e�I�	�E�LO�)��	?��|�rP�������Zˡ����-�)a���R5�˿*�MS��kA�/C)�R�%&�[܁���Q�"h����Wӽޯ�i�JF92KKG`���q�A�5�g�$�9�kc}�{���%�#	W]���
*��b���tF�-��^A(�N]0��Ζ5VKK�iee!M�i��'I��{k��:�[��U�T�H�5?��X���,i�lD��[Ց;��
bo�J#�(���ѣ��P��ĺab�%���q��i7�{���׶��b	�~>��)^R�BV���~F�k9���E�;�xJ���(1 ���׷̜_H(�43#���j�����ٓiya.����}y7�қW���?xk%f��c9�m+�&��A�˘�0�+��s@ԁ�[�r�& ۋSQ�a�
h��vuQ_�9��(��j^����2M� ������V�K����ö��B�A���>��С>
=Q�#4�ڝ�X�Η�<0�~��v�U�d�U���X�s��e�U> B�Mz��G����m���rT�� �%����AY��^K�·��N���N�Ǐ��)��P�Ov\��������4X�R�r+��Q�����$�嘮ٜD��B��f�5��˞�����g��D��Q)���~��/����"R�mm�}%�oC��NA�Vʣ����%�
��*�`��ѱ\&����"f��&'�{���<+��tҎܖ
v��>r,��fRh���}�/��>>~(�w�Fn���mj��=s[�.�K�SM�	����o
���RN��)
�D6�f�f6Y��M�z���U��=�Q�|�����5g.kg���%�Y������!c��
n�;��e�r�������0�|-�ū����Ѫ���)���M�X�aӊ�p#mk���+I��d$$�.�G��@l��m9+^�}�[�0[[f�1�W}W��g�5 ��A���R:<<�G o4��}����R[f2��U
M~��4a��1���{�n;��84�(��e@��U����J��e ���g�ۯ���056�7�Rv�Oӻ�۞���?�L�ެ�}���3���y���+�1����Mw�q�ҫ1�[(?� ?�[�G��HF2�{�n��G����"����R?�BΫY�Nw�J[W��,~+�h���%�:buQg�����VoX�(Q�W?���b�*��3����o/G�K�倄�c
�J��^�o�s8���q$�#��<�?^�A	S�cipX�rt�l�(�#��W��	*b��s�~���i��bs%�w-��tr|�6ַ�o��Τ$��$��^�O�ㅉ���RZ]^�?�pB:���u­ʭ���(�܏*�\�+C��al�vf�Y���Z��q�O�?8���İ���iv�L��|4{9���ߍF�R�Ȭ�}����de�B�E�`�i�
�\V�f� ±�,M8<���m $|?�>�����]�m��U�m�r�%cP`���>Lu�[��7hJ�*��y��+lqڣO�1�z���M�+��0��rs� ��U��̑�f�q��J�&��]~ݠActqw��v�%�qpj�8����r��8t_n``(Ol�z[^�Ki�sX�c��c)K{iCO�ۻ1sK�9Q�J��i;�6h)s��)�!PLb��ep�rx��*Չ�T�Wi\�����꒞�9�@j��+k�7�����7����2з�)A�V�@ӭ�����3��d�����#��@��g�KFx�Հ"��o����#��u'񺑙&����
G��fˠn
�8AGi3���
�
cŜu�}7����+����%o��l��`�п���^�ZO?��!�{_k3kˌmYg�yD>�](�R�-�p�_��� N'C3H{��}Y3"�~���F7��P�d�&����!���dh)+�Mg�غ?���qk~|g�(4��v��P�
���0�EЁ��f>(A����l�
�x0�	�j��٦�u�|���Շ����vdA��2eD�,�<pH{=�/Τ��!�����e^')�V�q��w�����C�0�h��I�c��o�����Y�V�Q�x���L�,���V&����L���VdZ�1Hʫ~�Z���e�XJ����B���_��(��k�{Uv7�έ�nm�Yɍ��zП&����;��B���~�����:BN���m(q���	r<����Ck�ON�<3ͺ[N�;�;K/��	���~������Y�u�n?�b4
m5�d�rr���1n䱣��3V��A$Xc���+)���Q�Ue{1���`����Y�p�!��>7�����&�N.݌�vAD��",����������H�QA�}������xZ�Wެ��HT��X�����9������r����N:�p�<�+%&ZQl����`�D�7xuq���j���[wv2(>��t��%��܎K3�(!��<�"��ތW��RlώY��t���WY4�n�f(P�U�w 0{g���p�~9Z�F9�d<��p/] ���� ����Y���Z[�A��S@����/��6��c�S���t !t����������oh�'MOƇ(�.�y>�P[�ƥK����7���O/ߧ����@u��?�G�����J`��/����w�e�(�c�A6��T� �፴�@��.x��ɠ�j[��h�Ӹo�࣑J���mt�عp���x;\&Q��1�r���ڄ��Ҳ_`�YQg��P���,id;W1�������5�'�,$�[�ijW�w4��XC����^=X����u��^.���G�aa�����ľ�l���`Q�|L��i::ܓ�yj%�;�H�YN�� Z�#��� Q҄ភ=��!kdzg�Wt�yb�u�?�����S�X��1��s��5��Y���i�N�=���*�?�ع��5�P�Ji��q����T֬���}�� ���U����C�b�� �P�ɩx[�2H���Y��d�3tl; ��R_�-��ix߂J�ZJy|b�%��$Na�����]fu#8/�x�����q�����n�h
� ��2?h�1Î��\����7F��C&����,�M�jP�ܦJ�-`�pks��P�-�w�:���F;�r�S�
E7nx�	���il�U����* �ݜn����y���~5n�I�)�g�?+t���=��t�{�;_���G��W�`dG��N�$+ȱe��e�����G�^ǡ��ӷwx�s�3�8�&~{U'`c`�r�i�"��UC�1��N�^0ʓ�*3L��v9���dξ�2Q8�&��A_����-n�x�&��/��e��� ��ݠ�W���(_Ьٵ����,���>�����x=��H�y]��>8����	>�i����8�p��pJ����0��$�� �>)iQ)ړ�	>;V�8�NK�3���_cN�Q1H���4I@��ww���~cУ�hXJ����N�ʬ�{��BI���g�d�W6�6��N��'�&��S-E���z��HGЎ�fEN��R^�O7�:��XNM0[ �	Ә��@܇��]w@�̫�c��6�|�n��#��R�4��x�5�^@�~à��A%���8|Dvҵ,��"!m0n�j$�W{���NjP|��=�v}�/�y�����c����<]��)�<����O�����4<��b�:���(��{	e��-Cq�u�0d[�؎Pa���Qn��L2�Za�N��A�ǵ�����%+�,C`��d��F9�p�N�_�"��\n�g���E�ӥ;�����Y��Q1{{�}B����'O"�Y��x	��5�؀�Nӳi|��[���9�<���/�m_���`����)M*��4�[��ilb�+�<N��;8��<��<�=�%�CA9�ɓV����	�S �yIYC�:?��vh���n��� ��n�p�B�����t9[¹pt���e�1sF�@k*
%M�9�ȅ�&�	9�*&�D�ͷ�1˨��������8��P�I@Qqw �*�ؖ�����E4��
OX�	Q@�p#�i"C�Ba�T��Ȅ�8䄣�ꆏ�F���uX�l���3��l��df�M�8�y("zh��g��+dm��\�"�x͇J{Rn�����))M ��<@�n�͈�>�fĬY����|g,����M��(3G��g�S�1���-Eh�Z��h��4�Zb��ĵ!wvh���8�����Xs{#�8<:!ő��� DC���(
�%R�']׀� �m������O٬�;w]�zyq޻��)��>\9K��|���=���� S��W�\��J(f�b`�L���M��^Dߋu�*{+(�#�P=)����Ϗ���tó4?=!�v%=~� -�ͧA��?y��s�ڧ͋�a� �o��s�M�Om�w�~I{�VbH�xP�<�5~r�l(��+ʝ�0cf7f�x "}��sE��(����k�pbJY�� �LZ�д�+Q�eX���s��̊�	̀_H�76.�
�n��L����sT�rۦ�r}SN��r���*�:햫���(�쀤2@F4S�;?�e��u�<�al��"�'�t.���Я�z��*~��<�`Zf���i^
�l�N���d�gl�U!2JdG8��>)����!iP�H���+;铔\+��FV����|8��̤��z��?����RJP�yE{�<䗋�2�R61�i= �ײY��� �m/}n`H��߳ʇ�'�u]4oXq:9�����y��R�W̧���44�r����Ƒ�s8¡S]ʻ��<+]��>����%z�
ٯ7�/o����x��؜>��g�o��PRng<���>x������OO���Ϭ�35����6�=�����І��b���,��3u�J_yZ���GQI��Q��c�P��|���yږ�������������ff��4�P/�Mj�]�G���&gTxO���ې��V����М���-o� ���ȏp��ti���Ʉ�B���%Lf�w��@���p�E�ލ�sZ@�+&o��J�D����O�_H���J]u#}��@�gnAGs�����*°�{�38X�������!>����Gr�,�mU` G.X�V�)^�tY��!�.،$a~s�4�	��3V@x.B?_��3��H�S��W��?��~�Me�#Z;�RL��C���|�P��@09��f6�߆H?�+���@�Vn�	�CN�fv�Y�]=�&�U��JO�%�4Hw9ߢ!��ſ����XF�%M<�y�Fe��@|L67;#>4�Y� lT�#��=mww,�I�`�lH���&C������؄�砑>�c��e�]��W���=?� t�ҼLc�������4��'�4��u�v�.5x���Mf�R�V 4P�-�o�yĈr+������M�p�rw�w@�u�L�X�&8ָGJG�|�qo�I�dBQ�A
:B)�5���E����㫄+��p23Cyo�k�����ysg�9�s����ڑ��tb��ckq+P���a6���)��B)U�5*W=�\_������#�Eց�/T�RxyE�]꿒79}_@g�1c��Zh�踅�s�C��,�)_�pt|�}�?|��G�,#�'��e�vfj�j=}�@J��`���Xf����_�?��4�b�1?�EVY|ѷą�+��	��S)Jܳ��vZ�����#C�SS�iuu�K)f���(��u@����f���A���*#=�6����Zv�AV�q������}��24v�A�`&|p�'�O�ťO�P,����~]Z0�=�D�nM��V��DVA6������)H<�g3�	���U:8:�A��ft�D` U|�133��'X��Ç�� �|��ے�Q�!{��ֽ!��
V"8aK�:��q9Lʁ�y/,Py�C�t*��x�������>��]�S���k+4��P&_�e��CN�s�"n��z%xa/�V��$�-�`�,C�s��pƍ�$�A:��
K�F��'ofz/ҙ�N���ӏ�{=*O�,�?8��@;K;;G^�t%!�o��tx������7Z(�
qB�7ʳj��2���j憧@5^�B}�B �}tl(MMO�ɜ��RnU^<�"�8�pG������Zӯ�2�λ�6[�i��a�U���Q_%�#�@���2s�s;�E����i�Ch��0�x��]o�s�M�U'J�ɫn��qA�>�5(�@����ygY�HZ�`���3��Ɂ�S	�aq��4��g����k���Iۻ���Ǔ���fz�n#m����4����gŖj.U^s��N�;׬�v�cTuC���d�Ca��f�P�N�v�8&�Z���g��jop�vGb1jG9�f�ͥ�?��]؄5�sߒP������k����^Jn�J�NɐO���}�AW���U��=�ӆ�I�̈Sz��^�aK^]����t���7��7��J�Q�~�)��P�"�BM@��\�`	U)�����v9��JŠ���z�޽[O�^}H>��59��>44�74�{��œ�P
.J/K8I��o�Ο�. զK~�B&J��(�x���2A��J[-|)�W�tz���&�����2�ݽ}���W����Yf;H!_X����i�1;�L��/
��dPNt��mޕ�h�Z\�!�7���cWD�/%���|j�K*�46��>.5f���a|��J+�P��/�Si#B����⭠��#�[�@]\^�c������AN��Y�O)c����88��� R�1*��\�&c�5��X�i�5�J����2����r�j�]���v;��l�ҭH��rc$�KA{�_M�2���h:�/W�t��n�&0���6�h-�KA�ca� W'���X��	e�ʌ����M	u�Ã#��*��ȴy��4�F�}q����(��-��֞��p�9�Z��N{��VEf���_�œ��BtI�U��D*�[�n��{kh�4�X qyP/U��k^ۥ�y���R�\?���VC'i�Ӧ7\?��F�v4#�D����ƶp�/�(Jne�iV�X@~�*�S4'f�N=�433����;�Ӽ�4����89�J['�����'�kyK���?NTs[���@᧽{YE�� *�w7�u�ff^�Ȳl��W�~�-e֧���q)�s3�iui6=y�&���:�Nh�(O��_��"�r]��{��.p�ם~�a�=h��Xe=��_
LTX�A}9|Qt=�J���_�ڡ����461�&��5���)�rc��ˋc)Y��oD�a9���d]>�!�D�*�~N##���V����:�A=������O����7��I�[�e��wE�C �>y��=^I�j�,��W�z/qA�Q�A! O�d��W�Aw�+P*��H��RX�&RI꫗Vny�F�bf�W>t���L�+siqi��Ju��$/谬����:�݀��"c���|�B[����+�y�W��`슃(Y�Cш����x�ׯ������e*��/b;�L\�G��.����i8
!E�v݀�ͭm�ݘ��m�����q����[�Q����dmo����렭�
TY��p�R9�����ů*�B�w٢����o�[�.�ȅO����"� �p��/uC.�Eí1;���DJ��ʨf��?�ȍR4���D�7�g^[LL�{fӝ����s=��?���^���IG�ʞײ1cgR>�d.��{y�-U����e)a|%?�3HЩ9umqa�
���*�P�-�{��c�⽖����l\�3ό7����^R�R�8TZ�v&���2~�@�2'7�ٕ�Eό�j�m]���,�:vs���Z�0L�l�J@��'c`���o��B	��Q�,X筁�Z4��?У��y���#c�i���̧%|� GF��!L��_o��O?�M��~J�Gʜ է��A
�
]2\tr)$��e�`�@e.%�v@J� J�����X���@Z^�N_�(���|�����!����>}��o%��h�i v�Ky�0�Oc��D�����@�5��+����(���;�dkӯ@I�s�	%�Ni��@um��r�%"=�<P�l	{��?z�@%���jz������r�[���[�]���t~�u��-k�h@.���L�~ĕ둮U�h��6���=�����~���t|t��6|<����n�ݝ�'�/<LK9����V�ʃ���2+�Jۙ�6m&�K�����᪋�	�B��5�ވG^�꫽R�C�eM�ֶ�۳Pn�brr8-�s�Â�,����V���("��� }Ml���zr5��}�E�d�g�5��w)>�BJ����>Ǭ��F�5��䦄��c�
<P�e�5��#vF����5��4(L�'�����F����Z��vc}#�k��9N�D�gm4���8[}"�h?^��x���哩!�C6��AK����]`Vj���np
[�~x3�0���zY@��zp���`�:��j a1�. Xw	pSe�L�rsT����.�=��᳓�@6��Ȑ�0`6�'��#u��S�3kq~&����@V�(Q7�L�.�̰��k�G��z�i=�OH���p��e֖u�r�@A2�V9�����d��7�\�]�DK�<V�'�F1�������gnYw����[�j�9�������+���Z�eD6��;!`"%��ܼ�=,A�u�B^�I������i�f�Ή���?��ܤ������Vz��S��~=mo�IH��H	P=ŖG�Iu_u�e�#j1�2s6 r�����H)D*�kf˘a:���]��_^�Iϟ����$�������4}��c�=L��G�9��&e�������vߊF��Z�q_���Z�	7�&�v��_wf�W���;e�kuգ�[O=5"�v%��/����o�������o�!k�KK����Y��7$�	%�{����(�۝�f����T�E��R8+��D�5�Lh�-��־L7�����X���=�B��MHa�}�y�?&���NXi#W����	Z�����+L���_����؂�+塾�5�7b�*[B�q;�� �'{�N����g�#̀�k|K_���O�pl �
�i:�߷Ó�[��,�b��6�Ax� �^/O`�2�o,NT��e��LKF��O�9�܁Aڃ��e�ă�I�.��;��ߓ9f�L�y�>���ޓ:���.&8~�����v�-r��X#�Y(�cc�2���󯠺���& �%�'���/�G�locz�L�4v�r�o�V��]>��\�L۫Z�P�Q5���_1(�Ɯ!�!
�+�qgC���V)ԈM�B��7D	4�=�� P�&''58H�]F		�&�D]�4��A��Z���C3��(��:2��q��/�Ց�� �u3�ހ�>:6f��������#�9���J��������U�?�p�|]���W���:��.�C��lb�/�(����mnn�3"C�/VJ���]=��3�gg�5f���4�fl��3]&+�g��J10a�8_#���ОH��T��Z�W�+��iyeA�k"KIW�t⵶W����������ͽt�A��Aٗ7>���l�4������A5�W�[h7�5�Ϩ�1f��m�ә�N����#E�H�c�z��M_�x����������GRj�ң����8�MC���B�Wʔ̳��do"n�7�j"�n�ޡj���*����um9�r\]���ݲ��w�{��������O�Y����ߦ����ҳ�Ӝ�Q���ɳ��5]��:k�cM7n9C�Iz9m�vW�n0R�e��vQ|��/�on��\]������Oo��/ߦM)���6��2����'O�<HOX�0=&I�Ti˴i�I[4�2��;2>v�7��0���+��a$-Jz�}�~�vZ�_��i��
9;��K�e��*��'���G���Bcc�K&��K�FV_я0�)))!4���9Jm�>�g���[����o,vw��Å����X�ev|ye�K,hG��)�t�W��z,���Ѐ��m���,��)�ۣ��z�6"'�l+SN�;�8pxp�e	�J�N)q&{�����i+�ղ�)�w�/�?#G��f��R�L�d���馽ܿ�Q�M� �4@��{�\��X�+Э�DD�-�UnTUzB:% 
M{g�N�e�K�fAت�ڣ̃heP���g���mP�щ�de��>�����JR ��qs1H���k)Q �O&�I[3��/Gj*���	�lKtDI٪���Yo;59jaˌ'�q�ת�ݤ�#)��[(!�ˆ�/�<C�F����d_AᱵjD�kDɉT���J(3�^����Q�Q٧��u�K���k��޻�]��A��%���-vh@�!��>�NHh)/��������O4�\y�Y��ե��8���tq����wFx�nG
�g�y��R`�͍gG��`��<�T�3B(�j���Lz��>�0��+��8c�ﱄ�e�c��|z���������~-��V�`�^N�c�
�B�����mvk��~����ԖY�e��㳠�u�/��[A�Xg�v��x8�c,�+W=�I!\LO�.��/���~�����Yz,E�[���蹏�'i"�G�,!�DY%���x�_���K��Ũ6��B�(�!KPNX���_�����fz�~�3��Ǭ��T�^�83ͱ����4'�k��=�9��P�s����=.�?Zy8@�����/n�R�T*hd<���gv7��2z�ޔ���6ɣ��(�Ef��v��V6)K_�	�������f/�?S���[��z/�=��U��X�o��A���a��7ML��ٱ��8mEwh9Di�hw44
;������\�6�6���k0�x�.fm�A�Oh��b�`���� �m$�F9fxܳ���v�1��@��
�i���^�	�fv���%� �{���t�ʐI�k@�c,������XC��S"M��w\w8P�Y@�{��B�����3���L4�i�`.{:U�SP�����7�(��E��'U^I���8�jjj�3�<a��t��su)�(�.	�CC�'�.���n��ԇ�<#l�{'�>��Rf�7Qª�1�b���v)��z��N
���&�A�=8�J{�2/�v��]هQR���Wŧy���h҃�
����,Y<���A��UV8Cq#k
y��(�<q�k�a����FJ�Iz�fͧ�,ۗ���!�A}�x� �ĺܝ]rɗI"��X��@	Ӥ���vd���UB�(������4'�����?Y�y� 23DFDj]Y�X$�d7gf��<[��a�����孭��ggzf{ZPK���Ef���uw�7"3��M>��s���p({�����ץ�s֤���=x������L���V�?�෴*����c���o`���9e�7FQ�ƞ?�P/@u��Q�f�rV�X���Ͼh�������S&x}m�Ň�i�n���X��=q���DгҀ����G�����肕���
X�#ANYU��i���E���͜�����_��'�/���!�ggU�O��0NP�9�Ί��7)���B��?9������o����:�;��%��߶W<�A��r�ӣǏ��E'���!��ĺ�����kRp5Ѻy�_Z<'Y�Z����G��cX������S�Ìe��{˖{��-�\�d5�"�W�@����K_� :O�XD��K��c9L�K����BF_���T&�/�q�߈�0@'AVD�,ɿ�=����q.��-q��y�W�>}�����={u�ԙ�U_�/3Bv��_	ʓ�:�Ѐ9�t��Qmd��!�〤�1"��h���2��Ę���4�xR	/����}I�;_�����%@�)�F�&�&��	���Ϙ~��6�{��#�=3�6g���	`y��>�/�R��>�C7%��>b��Z���QI��q�鞁:Fa�ORX|o0��������,���<��^f�Qr�T9�Pzа���ʌ�ʭ�Pnc����|gw?��e$c�4��RV����Re�=���U��4(Su�����ZÞ���+�ӆ:���"��T�}�UebW�ہ�+VQ��ɼe�gY�<��SpTh�t��a���߄?�1�1(s4�]RX���TN�ߏ�"�c��RN�Y}VRN�����?H�S�i�,s�����5��xA�P�>��sS�+m�º�
9?���?x����o��_�o/���3YQ=<�b�I�G?qW���?����S��\:�����Y���2��}�>޹}���G�a���.�d�$��"
�w0�0@v��� �Aظ�~�Y��U�.��]d�]9a�e.���Ǉ,�Է8꩏	��U�-TLB��)�*�݄��>�Ӿ��G2?��t|����I9�^m����Z�4�m���N���Y�fDwu�ė��L�=daXm�V.�`�4Vo}���7�x��¸f�o���K������3�Ǩ����WiM<F;��0D��+�}����_�T��S�|e�q{��I��xIB!hG,(\��������J�U;�S^xD.�Ɨ������<�n���r�;��0���/�ޜU���vK�=���%���kk�X�I�VnS�s|���CIm!��9�L��[A�O9�应᪽�o����+���#�n9_7?��H��� (*2�p]���2�i��=��� ��s��p>J��������lP�)�?��,I�dz���rp�r��at�K��CtX��wW�@�E�˲b����t|��Pn�\�$EJ��Z7m����_XE`s��*�WK� �o�J�T��s�ҎA'g�n�r�|��^�ΟSX���x9)U�U�jϼWu�{��hX�C�OF�7�ɾQ��Z�غ 
;Lv���b �3�gc��ω��ΖA��8��l=�bˋX|���V�E-�*����G?E�1�ʁ��f�@&�{�Xё��	 +�t��sy��u�P��_��Okۻ|�n�ݓB��?~ݾ��;�C��wL��)�,��zm�
br�^��m�����2؎{`إ�
� ��.K�����ûwڇ~����Y�V:�ӧR�8ll�?����7��|���R��d�4a;(�u�{��AF3��}G;�Yt;���V���6<	HS	�����J��+N�ˌG���g�������s���>��-I�+*��K*�K��n��?��}��?���ޢ���x(%̫��������Q
g�{�U����bXʁ�R�:�c�7&�l)�S���]m���m�i)t�ڕ�������[��g��\)۪�T�8EBi;Y� tJe&�{�Q���� ̨����ҵ���������Ĉv�C�~Zv�]����˚��yg{˲�rB[!�w��D^���_R�	��+Kc�Q�+��K���6�zks׊���2J;4y�^
.Os8?Z�9Τ�����aO ��9!Yt�O��a� b�|+}�9)�(�O�rs�G���$Y�XUG|�G���5���^v=�~�`��{H7RM @����t
�a>�"8����ꑭ��:uB-���@��J(�"��R0�7�)�dR�{I	1����;��(��m���[�t��t����v�ɡ �*`�G��'˟�z���'f�+8��Bf�d`E���#���S�,�8F9�8ޘ���PtV�ȗ� �"Ù|�y��щʢ����(7![oD̼I_&�[PQ�x�
a9�U?������<��ԕ:e�9��2�H��p ;7���� �M$���G�t���������4+]�������K�OڣGOU�r?�>�pV�#�ŀ
�_�C��2�|��U��etT�1*�N`�����UՑ+�.�;�n����~�n^��`��'�7$�����7��W�g�|W�G�u��G��*y�-����fϷ��z�	��;��:���gt|��w�w�L��}aq|X���񿿼�"��zu���x���}����Nu������'G^�Xi7�]jw?�%��n޸�����|~�5o�[�$iV�*�6*W!1h���P�0(��1i��(�B��-�,��������6���3GH�P[�?�ԔR黡'>�^P�b�FT13���A p�7��7�\O�$
�q�����#>k��G)���"k<����$�OM�l���`_�a���@}�y1p��`���Ѭ�=6U�,��-Ug�ǂ���m���I⺞H���GPp���(�E��<�b����8��U����?�؞��[P}2{m�>}�:��eU{oyO���#�@��6�r則�[h����Zir�C�Ⱦ��vPN(�S1�~�;f��d��1u?���
�wZ4₨���%�ܣ(��C?���N����)u���j����<�G7�;�j���c��Y���a����Z)�6:�h�����/b�2�I�H��Ș�[���i~�	��B��&5�A�A-�j���i����,����.� G,�#^lP
�o�r���;75��h�<��W<"g������ً���x*�W����EY!�H�ҏ�� �S��
���b`�2.�t�<�Ce��cl�`�8�c�, ��ύ�(����r
�[��=D�E�J�|��R&���u��^+�(��jKI����;�o��>��}���Rn�H�������W�4��z�~�o�W_�����*�W�,�@ز�����nd4��U���\�ʅ��[i.D���{���C��#��	�����N`2���	O�έ������u�u�mm�o�~�����4y֞?c�K����j�u�M��	͝�w�>i}~�2�g��$�����ww@��O�\�'�T�c��!�+	����֎�+�qrܟ�M �6�����w|V��/�R�y�W�7�0����\��O���ǖ�m^���#M�>M���®��k��?P���i�\Y���������1�a�y��3�P��G�l�@�];�*��#%7N��s����@��]�Eq㽂�!����_%&f��&��ڲC���~p����D�@���i�c�B�Y��@���y:�Ʉ=�B�H��M?��ݻw�g����C ����~��-�>L�<n��D?��QiP��H�n(��2��@-����.�|���|/pv(/���|�9-�@���#0f�}3���b8)��~�
�.����6�F�)	�@���\;/T��E�|�ȋ�we�w�š��+�i~���P�*��tQ�\1��II�a�8\�X���mDi�#ɋ{��^����[y�M��<���֭���s�C�B�B�E��\�����tP�듻��`�׻8���}ٯ��E�����V"��B@�t��cd(�7�},r��?,d�f+{9O�/�1��;g�|w���}��ѣ�L�`���V'@�=����ƛ�(�h�!����L��h�����xe�����O8���Rp4�sV��?��iۿ��OV�8ig�U(=:/]n(����̅�-��r0����S����� ��;���l���Gu�qu���E �N�x5�1p>��m@����ɤ%C�XI���B�����j��ӄ�ޓ����d��|ŏ��(�U�}W.���7��Ų�?����W����=)���z����4�άH��s���Nev�����C}�U@&��!z�8��9��ѣg�Oi3���@T�&\V�e���/��2	�p=�W�u����J����s���ӊ-�Pn�}���L^����#�|+��+��s�gݢ�}^^"ϒg�GJ�����ˎC���4����r21%��[�[y�bȏI:�!_�w�ܪ�0)�r�CP|'X�K��,���ʇ-�}�p/�H�Q/��yۚ&FO�>��N;�lq�e���}�qP):��fӐi �`3�7��2��kp+<���N�Ơ�[�nׅv���
�OX����B9�����a���E��@�8L�C��ʴ�����n�cb�����|�;�Q�i&��Q�ܥ<�_�Ӕ�a|Ί	����2Cg���֞�}w�(N�'R$\!��0���v�����JQ�@���;�-�K�*���#�z��A,G���]�垀���-����7�V�3��q'�m�����>t[�)��k�>���rʃʆ�ærY��.Ō���`I�:��?�Nn\Qͱ1|�
o9kpF�}u��^H��4��r�#=�9�
�x��~-�p/��z�$εյu���JH���	#�Pn� ��<Ņ2��-��+�/��E�v���Z���+�Z��Gw}\���dU��{�=y��~/�������?��ߵ?�鞔��9��EN�$,�p��pu>�B�O�)�����2���r ��(���G;i������0x(��&}L�LFS�Y!�����=�}ߴn�<u�2YZ���x��c�?}�m��o�����o�#MR����fg�ō3������'�ۗ_|�=�w�\S�U?�ˑ��>;e�id��JD����q��O (�(�Xu[n�ޜ�x/4q}�󷷽O�6OP񯭞�b��>�}]��5)_q���+����$R�.OX�*��7#&�ϴ�I��ׯ��Ӧ��C|�P�bQ�	ߥ˼T��{YJ��&N��Ԅ�V�*/e���z@�cܒ�F	!N6�.�8���2a����m��#�X�G�E���N���s�ӯ5�Ef�-�ϓ�ն
f���(���-LD4#'�#^9��Q7{4Y"_�۶��-�tH_�ME�#|鎗���&�]&��-x����̨̅����-~ƀ���k!̤#8!�,�%�H����<�,t]OYT�S�f�? κ]a�!N_C�S�f�b�ߜwyV|����ɥ��I���=y��nG@x� e(WF,��I#�q�a{%w�%V�dI����<�p��g�]jW�^����4pV��y�.�p�;_{�62e����,��}f��C�NT.�1T��ϽQq��#vu8��*/]�+y
$X����j��n/��O���[���>a�D�,{2�w�:�ʷ����P�)������<����lb��(j�{����ۙs+Rl7�s�7����ѪLk��0d�u�?��$ϔg��p����oⲗ�=�5�$
ᓧ��ᣗ^�dՇ�Y| 9����ʂ�	J��Pv�θn $�t� �F�dd�  y�ˏ��"��5/�쩃ծ\Zk����nI�����K���V����Wl�o�}��|H�QB���/��W�Ӵ]����[G� s(y��+pP�qH�	ԁB�{�E#�����%=h%�b3�_�-ӵN�hwi��C�t*#4J����K>��:O��[ZQ�9'e��O8��w���}���.�=)(V^4�_���nߺ�>��z���|���.I!8�n��[��yK���੝��ު�yP��H~�V��A���o�}���Q��I(�~Q�����C��K��Ź%����r��,_-��Y��}�O��G�=�AM��i�����k��6�r�-G��3J���]���1/�j� E�7�)>���������.���6�0��C&��� C0�݂�(���e�E���({U��%J����K��I{�䙕\V=	�D��9v^<Ռ��š��ê�Uw����M��	":�Nɋ�;���4�V<E���,�D��=�-�͞bN�9�lS�59M�YQg�����"m���z�2����!����P�B��4{���������@@���,�mt��o~ұ� 画�%'��|�\9YyO��D �"i\�S��Be!�4h��,.�# q�X(. nUY�qcS6,��T�^~�uuP�i?�f���;�~��MP��8�y�S13{��Rl5ڜC��FJ���#u@oڥ��ۇ� �޽�·O��@vvx�t�8������~4��nU�|!G��?�̎b����<G�� �EO����$ڟ�@b�Ȭ�]�f�*����u`ey��
�UFQ�|��M���3�����ַ�5^�K5��[�>��"9�lT��t~ɣ/��~F�?S�ZX��|��@�y�2��pWr����c�8�+�k���?E;�����K������bs��]Yo����zpq�gx{�R��(�6&��5:d�0������0��A�|�_<��HRh���e��v��F������?�����O�ō�e+J8/��{�mnr:�0uI9׀�
��Z+elq��ʚ�wG#^]��J�F�g��K��%�MMn8�wiUyQ]���8δݖ�r$��sOo��?�Ţ��d��̞?�m���ߵ��_���韾j��=U�U�ZY3}q5��e�$0�3na��'�u�A�Ou݈��8���a��cnʋe���yE��
*��B�8+ܐ��A
��p&~@���<���OX�.�Mf�`D�P7�>@#&��U���y�����${V����&(_���?x[	/�Vڼ���v��Z�����ﴻw.���-�l;�O�k�K��v=��I���u��9��]Ot�ُ0�T}�P�=�7��(���ų�c���-)%��{�~�ǯ�����Ǉ�p�/���W��~��-��=1�|iC�����Q{�/�A��X�YJ}(Y�,����'y=)�g��ҹu������@�o�=iO�fv�I�_�Z�Xj׮��5q���kmC�.}O{|�,�'p]A�vJ������]o;���F�-g����D�@?L;�q��'/�ak��~������i�������
�U��W9'��]=�.�'Z�X4�J[ħ�0�_����Vl	)��� i��T��7�'퓾�v�?� �[�����7�f�9\�o
���ۜxBf M�e��p�%O�8�<cB�?�q۰�R(B�+2�B˄�^��~�] ��Y��]0��K��t�cͳ �7�'���>@莜ˍ�AM�MX8�y�ԕ�L�%P4�A�{�T�
4�ԩ;��#ABt�����[����y��t��k3�\�ؖ,���NjU�qd��қ��Nt�]�쟽[�)�f{~����U77��F�tV�T�kE�ŔW��aA᫢�;�f��]N&��Mv��I��-�C��-�%�P4��������g�9,]��q�IE:�6�H�<:�8��0S��2#.�
�o��S}}��t�p ���ͬy����3�]Q�=l|۝��Μ�R��AR�ZlP��c�-���t��d���DvttQ����ɑWA�4�忾��|L�iqR+�L&��^�/�ۣ���)䬘��R<1��!&L9Xȓͦ�z����OL��|G=Ef8ś�tP��w�VW�x/�����cY�
9{�xL	����~�����~���?�P���_N3��0q���*!���!��yIp\L�C���+Ȝ�<���7���(�I0�5K%����(��9�̴
�����Uv�		���$�*���9'�Y?�a�����z�o�{ڞ=��ct�X	]nܾ$E�J�#�ڕ�RjX`[�&���1+�k��Bs$,����ЦP�Q�P��������˜��KZ��lݿ�Pm�&�V��R�y�7�s.�MҮ���t�J�b���?�}�
�����0�W�-����+E����R{�b�_+{�bS�d��ϵ�g��V۝;W���՗�� ��\���.��ng�~_ծbb.뜿1�,����4��5i6NpI�'���5O��	�`����o�)����ď�"��H��`��$�$O�⽌I��0�1����㍟�i���:L&h꾼�����,�Ӫ'-OL�I��r�6:[;��7��0!����A8ʘ���٠`�۔�,�	2�(3Kƶ��'��0R�n$bV����R��1/�I$�J �_�35虐�!Qa#|5��� w�a5
��t��9���zJ��� J�:Mp��1�
�z�A�e_��x����ڃ�G�s�o��\[���1���?w�Y�gr�Ef5wD%�GKL���T�5�-�H��Ov�%)1�YUdV[+�$��?��U=l�x	�����3|������#ٰ��Ǒ��3��W����Œ7b���Um�汝��e)��m�o��7�/�H9$(ꯎ��ȖA��2 ySV3�U!e������s�u�rwم���sE>�Dv(�#oia{����2�������<�����>���7�f��\������=��4��d � e��%y�Btx�Y������Dn�ݽ{�}��Rhn�W��f�
_O;l�~�������_��3�V7b��W�0�nw�C�g����s�� #& kV���mM��(�<v���85A.�@O'��r���1�,[ɾ�kn1@N����E/?�W�o��;��n�0~H7���쥶��9�o��կ�~�����k��C�K '�x�~��&:�R�P[�6<ic!�UQ?a�~VxT�j�Yi�}1�9��3����D�z���������˘>{��=��)����O��I�UM&iۤ��@Vca�����¸��S��Pt��-��P
�?{!sS�:j�"�����s�q󪏚\[gO4�K&�@Q����p��)\ �G�5��lP y�y�G�/]�m�ƱfK��/'/�=z�VJ#E�N���&���.b^�9#� �D�6�׿�����Um	�����YH�P�������Qn��ءm��@�����I	P�m�iWN�Rr��a�u?�u�� υ�c�9#��ȥ�u׌�'����py��b�B������ퟁ~$8s@ ��Lb!�����HT��p���g�&@*iV�c����E�.a��7u8�g��&�T������NrU���V~��Y���RD8"eooO�:PJlB���L�c�s��FC6]v���NPf�t��ь\�콚R��S�����t�� ����"o`��'Oۖ:c�@`�/x�qD��J,�����"��#Ԣp��ڊ�l���ϻ�i]�rُ�
�ɽ���'#��?��\ؐ/d�-�wyf��= &��O4���� (R���I���loa��vC���������ŋ��������<Vc�";��`�����t�y���Tg�c%�[^z;w�u۸��-����}x���+��Qlw�^K��m_}�H�Ͻ��7۳'/�K�g�g��z2�� e/�j�U��Cd��9��|G<OhUQ�U'C���� ��Y��z	Ԋ���z?γ;@����V�!�=���)D��D�zuۧ#(���Fځ�{@��>I����񓨇�����[��LnՎX�C��o������On���hW�_T�V����v�
��RdX�0X�^*��c!�,��%9��m�2��G��?z򢽐�˩
�z���8����K>��o��t'y�`��nI?ܗ�̲!/<�g��s��������ec�?ū��syW5i�"�b�!�s�En?���IU%V9U�<�g%޽����8©/��q�~�ϳӯ��JD��Af-���i�$� 3@�y����b��M�n��[%� �������	cR��¬J�=���Sx#i?�E�닁4�t�����l���/�t�p?ID����gȍe��N0���C��l��P��	y;�s���Z�Nl�~?0㪐�J�Ĭ�\��6�Iu�
@R�l���Kٛe�|*�պ��a�k��,p�-�[�Ͷ�����|�!�`�;kw؉yｑ��ŧ�W���p��|��Y���ӯ��h�چ:RV/�C��ض���,�j˓�O�3���f��&�<p_o�6���\F�	��8k4u(<�#QxD��|�[����uϮ����9���6�Ӛ��*U�=�3K���
>��EH�.��7�ó�[ɛc�.k ��Rn9�k�7E�����H<���ݿw�=}�T�,%a'd�ƴ���d��bC��]
�(�꠴�X�=�*�����ڗ_~��܉�𙰱����Q���^����u{t���@f�~�G1gd�s���e�BJP�-�!���"x8x5/���ա��@y*|*j�4a�˃
{
X�����d� bԪ��{�/K�ݓ�k)
�����m(8+� O��3�����/ѫ����M�6U�X���$��%o%Y�-'[�O_���_y�ɟ����y`�yt��wۗ?�����O���_�s�l�!?�Ӭy�%�B��N�'���$^2	������d��d���I�s)�l��T�s�͕k���_V��cd+��!�)�K�U�����%�ݎ��H�'_|(�OR�r֎�;��ҢO�x�b�˗L�y���#2��4O����(sF���m`>���nQ_Pnyѐ���Ix�[>HsE��׮���.Y!���"�L�X�o!ς�$�n��;�����ezզ�7�w�>!�v��}��w|.1c�(����?��d�W=��}F<����i���'Qϲ^ͣa����>�Y��2
 G=�mb8��F}�26)��t�g�if�0$bL���b�����6����0Ͽ�4[�Xy�\a���+��+�rC��HVl��v������#��Ґ.ng��B� ��#CŁ�Q� ����W���R���~UͶ/k���X	�w��Q�ϟ��b��Oxz \Y��3)��s�5�,8�	��M��hB�]j��{���v�r|��H�p�-�?�"���żZM$,r��+�{ݧyz��� ��"D>��U�blG����T�+�/�_�4�������с�����x�<^z�����b�TA��<2H}Ct<ᆖ�b˓�˗/�;�l�}�q����x�h;^<��9l��Y`^.y��V�dM��������b���� ?�'��Z�-7�! �w~���9�b8W�'R���Um�-@&�,����{�D�8T��z�	P~���m[ᢝ�K�e�V�VT��*�0��(�Pb����P���m�EQi�ڵ��}��?}}���o��~��_�c��X؞u�ƥ��'��O~�I�D�.o�S�9��8M�� H� �ŀ\�oB�δ��(����>B�������^��G���\��DX���#xM�ŎC��+|�:
�v7b�����G�o�~�e����dQJ���?
!��<��[&��'8�t�?a`a!��e��c�-O"�n�r{�UhV8%&�KN�X�c�WnW�3�(4!ꭑr3�LL������Bś�g�±M�dQ(;e��cW���m����/�-k⇂�#/p�/�;c� �bP_�n��6c���[p5��������e�����5B�𶄘)T�y
�w����S,������S�{Ht���<���a�< �:�y��e�K8V!�?�}7�� ��>N����*��[^�|��`����� _�h��{�\H\:Jt؎��+��YQPji�G�u_>�����v�
��X�eu�����	|��Y-�8v������ތ\O�a��m9O�Q�UF��;To9�]�p�mll����7R�,>~�O����҈�ˆ�3�*_	6�~:�9��h��M.>s�> �CxeTi�:'��/,1�sV��8^�tQ����$������s�K9H��m��)��yp�!�!݀A:�Q�R��c`�*��Nr/��\Q8�ǣwn_o�~����[�۲[^��;`�v�J�7_?�l5qP�X^]kkX��q/+���=_Zb�� .�G\�b/}���!��<��S���V4�1��&�i��Aʏ�q8	Y�C����1��T�sh�h�L4��,i��F0Y'���R�p�T�A��]�u$��z��O���[�%� ��>|����?�����]�������؞����ƹv���嗟�/~�&m�g�_@)��+`���@��쬸UOq7���=�)�*s!�%�z��{�����Ylp��~��{|,�_Ӻ��'�D'맕[!�T:1��{�`?3i�������� ���(>_�gxy1���<?T�A��[��ҿ�_s2ʢ�	D
��i��u��b2�.9��cxw'&TVn��}.���|�����r�8�$�҇!��s��r�.��x#�=̼)@|E���X�UE�<֊tma���g��b���	�i,dQ>}Rz
Dm.��0��98���(N���\%���r�m�Ӳ=B��h�\a�� &�=��f�*�f���H��Ёa��>�M{��3�}�iF��!�m8��!킻~�K�����N���6X��Qc�=ǉ��������=��e'Y#rI��vW��������Ѝ1�q?�;���`�+i��@�?!�4\>~@�������Ϸ�$���]��j�E�0���7�g���p�D`���Y:>\��:P�e�e2>B���Ha|�c���/¡��*�Q��E��*�Z�	 (s"6ʖ��R�4Ƕ�P�Z�Z���l1��ז-Lx���u�mH�}��<+��ӊx�WJ��K��a����g��J�;�ߡ�s�8����>���_"㓠|��:o>79�a���wR 8I���(�^�I���,��������rÀ��:�\YǄ�tx��-&��O�Gip����`�f����@�(yh'e��"+e�@Ȏ��	��{�Ҩ{嫷7B+�ԙ���u��/H^�?,��6-^��$��\�p�Ž�O�������sqٞ����t�?�p��Eݳ"�t_3!���L#US?	����"T��L|����c���rN�����E�-�Q�P���:�^����n����1�|��L?�e�'�\��eW;M���g���Pp�3�9c�2#���ί���SJ��
y�S1����4�%��Z+��	��l�{Y�e�����k��x��Z4����%s�a�½Rt���U������8�[}�ț�,�GۄO���3
5�c�������KK�S �8�n:��xuJ�������'�0��Y�4����,�� C�ȑ�?�Gg���`tŬ��";W�J8i,ʽ r�CJ�si�W4�e�T��Cez�(#�J����JI�e��Êj<?H�����t�����fUMۘ����U
<)e� �VF7�D�10e<p��&�|[Ⓛ��	F}
��]�Q����"������sv�
��/����yL'!x���"��Ŷ_.i<�ϯ����V"B�$ ��y��&t ������HSb���j�H7x�O�*l/��h@��� �b�=��}��D���o�g� �H=8"#��20G�Q��.b*��e��,T���ƪ-�=���2�GVp���9)�<�{���?}�#�>}��U�x�=�K�fR`VB��<Ə�'�F��W�E*Ȑ��s�����@u�� ��/�O?��}����~`:xe�o�{־���KF�[���)����� j3�D�%��˲I~̓�Vٍ�-�	�2+Ң�\��}��ز�=���躧(�]��R"Ar C#mK��K��=d�"�sO.��'軍f[�nV{��ґ&����=�շ4^t�d�}�R$�/)�� ���o�!y*U%��S�T8���j�Y�tU%���
�>�j�}�7�7���	$�X��$�KW�M���s�툳��8��%���Yn�IVx!�B�0�����;��+*w^,;Ҥk�=y�՞?�F�w�\�/i]���~OmpcU�^
�~�Eu��gO���+�@~�!�$�?L��3���gl��KL�Tƺ��^v�����q�r�뢎�W����Bg��9�k$�L��Nɣd3$}*��f�4�Q@�5>�i�L����7�M��E5<'�>�~$��r&��eJ���ٸ��@iV ���0�鹭�u�	,�w�3�q��f�|��R�(K�!�������}�C"Ϥ��Ѥ�
����8r l�)Zl��n���٧�#����dD8LYL�4�>������a�i�S��W�Lǂ�����>P���@� L��'3$9���/<����ᰎ��[��g@4��$�C9��5�����@�|e�=2mtA����k�7�����K4�dz����e?t�N�i8#��M*�X9+���4q�ZL؋��ø4�g����U��pv//Y��5E/�D������o�stvIAt�E):{[?
��s�i��) ܜ����@�����[�BV	 �U�&'�?���]l;�e%`*�(�X����t��ǒ(�LHVkѴ9<�-	�������K"�F7[?Pj�	ᙣi�/��+�1�H��5�$��DR

2`��u_u��x�x�k�;7����4��JAeGrD���)���Jq�R�`����d�v��-C%}������	3b�����>R�Yr��S�x��޾���0�w��-9�=(́�82���[�&��?u !?!�����#��]Տm�-�Z��i��Q2�J�1��lG���4"{�#L#\i](��xKm�OVJ�c��/�� �V�uW
/Q���Ϸ۷��[�?�X0)�^��~�x00��}A�;��+���xe;@y�r�mnx��f�����R��z�	��?�gV��Q����Ț�I���6S���Q�a�ې(o����=+�<$oj�^��(-�޲�2u�dȟ)&�Ѐ�aQ��!��@��ø�[�(��N�S�	6���"S�!��U���}l�P���>"�8�[����)��r��d:�8�M�;c��=S=�a�ܘ�������
������ �L��L�ۈ���IF�q2��P.oÞ�z\�x��E��&�%`��(#��2�y)p����Z���PI))������ 39d�y��C��*��S�-�����Wt	��Ȋ����:�u7�R��B��Gb�+ş����FU�i�i��o�#l:�݃G�u˵h:C�R�b�~�8��E:T���oWZ��KgO^�r�U9�Z��Wi�ˡh�C�k{�}7 �b���8%���k˛ża��]��=���E���!~�3���V=�a�7�*Cp�(V�P�B�eՑ����C�v�E�uK���o��ޖߠޔy���UP���*	�|�Y<��v�O��W��
�ҜV-�7|~T���������뗥���I	�C��Ko���@�ͷڟ����=�-��W�̋�3F}4f�Y�ƚC���,�V������5��g�y_
��&N'���煮Q~C��g��bK�(�9 � ���3/y};�M��+Vsb�(9�Nx�-�m��	�vǊ���˶��*�)D���./𽔂�����ʨ��2�IQ>š̩CN3�u�u�L��xu�aē�{#>�Xq\O���ч����n�]�=���R×��#_o�������K�8s���E�M��,�Q��x��V��&�L�&�6�*^WT���`/��q�&����T����ۜ��S}RVG�QNS;�\b@�k�'f{ݛG��ٓk�����,��z[��(�
�&�L~ϟge�j�d�^|��z��<&n{w}4,�E��<��4
u��\�n���l�d�ef�/L�>cA�����
c� z�5_��+DX��D�1����Au_����_:8c'�>�u���ΉM�=�'�?�Y.Se.���`����|;�c�q���T�0�	�B�6��t�D\9(�"� �O� ��Ϝ����(�S�3�� �sB���Z�	ĪĲ�k�+%T~^�W����ǅ�`EK!�F0�{hX_N���6�wf�^��L���ŀe�y��7)]Vj9~&V��:"\ʌ:[�h�1�A���QU�*]�γ��8 a�pҽ�HX�3��#���\|窔[+��$����m��;_��z�/%7'Q���Fv�W$N0���7d9+�!c1��ڲ��B�ɋ,ׯ�,H��.�����/�j�^<�q^ދ�0�����=�p�ܠ��
Y�΄�(��^��^�;w����hW.s,+9���m�Ԗ�G�;!+͜�ţqȒohF�)������X�� *��e����O��<@Vq�#"(�
�X�`����`ޣ��JSz~/�2�n�$DK�b�O"c���mK� �gY/]>߮\]3^�9���:��,LPP��wLb@A+�yo>��c��x�?V.}Ԗ���9G�I�3�(���J�Q푽�W��r,��89A�cLHJ1#x\�hL�ȓo�R4ov�$ ����<�=���"�:�v*����g�4i@q�9����Mq���~��_�>�Q��X	��l:��'�й	��� �"�X퓋�%�K��55�,��?�[��-�����[O��#t����Pc�]���'F���#�[�4�%/�mg�P�����/]l�3����۴Ő�IPIv�	�1ı	�.�z+�ծE���<  ��IDATM?�Z?����;4<Q�T�.�Lκ]���\d2�e�O������P����p,��c��y@�`�� QN�6zV�s 3ѓ��+��d�͗3oo�ol����f���&��ܪ\�嶀s`Ql����6����C�%6t�+n���#�����_�b�OG��2�*�M�¼�{�-�e�>K�uy�#Nx\�j�38|���ܲ�2����!���F�<!�/���G0��y�N;0�
�Sj�m�����+W��K�5�f�D��:^������^��o�@�Լ��L+o'^���TiLy"���^N��-[?�69D`п���ʭ���S��AlIx���ﲢ��Q�����)k@�V�d-&�a�^�v@�f��U��8�Co�0ݸq�}��m�y��Yq�Z���ɓ�v�/�=i�=�1Q�
碲��⳽1�QG\O���.�%�P�,B��c"�^۳K��D_CQ���~]�!��<�S=������v�ٮ��� ⸮);n?(�NԮX���Y~ �.�/�	��s�������7�?����o�~�럵�����O>l�n]򙲔��Go� ��#�J״ �Ө��(�`�,��a�`G�c�6����r��}��ۮ&��R�Xq6���&HL����Չm%��8`�?�1�-����V�(#��|��㣄�O���x�m|]��Um��1&�7�&oݺ!�e��3�HJ�hTO����$�1�eX���C_�z/w�d��ǁI���[�~���Ue��-� N��2�:R�P���!P�TNB`�@��-O�|�awg���1���"cx�y��/'�\���r�ϝ�S���X��m�U��,��SE@V��J���Xʆ�n9ޓ�O(�%uq�j����E1�eI^���#�� ���r�<*>z����\��?c8�.W�Nb�'�=	��T��?��	)�Y�Q<��Bpn��B�#��:�o�?�	�0}�j�,����+�FU�c��e��ݶ�����b[�i#����8g��01̸p���3��ާ�A=�~N����ٟ�\tB�+(�4��u�Z��u�
�TzE�Wq��D곀?!�p�v�=A$(�Rd��!�!���H�8�UZ�1�b˧$�*����=�<mU��"��p��0����4t�}::�)#{CQn5���۷�����=�s�r6'_�C��i^���(��8�Bt��d�6+�! �rM����)<R�E� @�������Չ��V^.|�t�=x���Y	c /g*U���pDKÅܤ�x@O�ra�	dА<��3BLbx��[�D�y$�H�\�+y]|ޒ,o޾֮I�/m+\(Q(�G|� T�� f\1hK��~��\����Q�T5��N����%G�S�7�ܐ�/�I�ۿ�i�7������~�~�o�~�7��>��|�x�6�[5�_+Qb�V��~-[~p�zjH7n�Ľ���M�-���8�������w��[o�3��n�"z��uO�xq��H��x$[��Y4r�ڟ�>�P_��w���O��>yY��^n�i)<�g�v���vC<��>W��c��Yn������P�Բ�wTl�',�w��t��&�a���F���-���zݏ��H�E��k[aaF�g(p��Ìk2�=�e�6��r�w΅E�$~��rޭ�T��<��~B��l+�D=m�`w����@�#&��
�y��Nt��rK^���nmkL�c;���,��wʣ�lGY�ݦo�0!a��A�]um�������.�fch��O����e��EQ�y0:� �(��<&��A������L3�+��TRc��]������+D!��EPA���#l�u�Z8/�.��B�B�B��[٬*�ᗮ��i�|q�>���Y��iUBB�WT��O?�w��K<�ݸ������1�g%�H��K���&y`�?����0��UW��J�4`�<�c/�:Z�����u%Evyu��o���{�<#�`%D�!��)�T�qW�����c�ߗ���y���c~��u(w�m�i$]d���$yEB��B9��~�c�w�#j�甄%�v�����C� Ճǧ���G�<{�έ��յu���z�%�
F��4�(:tGՏЪR��Y�Gz��J�eܼ�qNW�M�Kj 8�y>y"���K)6�mO�.�ٍ�.P��i�\��8����,T�<�4�B��b�$�������G7ڗ?����o*�Y���>o~|G�����x���4�4��HI���_Pu�ړ\��-0d�1XQ��_@����J���ͤ�{Z��j�F�\��>��n�����������?��_���~��ÿ�U�;)��}z�]�~A��$��c��x�_��˻��`��u~�n&����ogۉ'޼��z��:�ݻ����oۃ{�����ʊ']�=AJ��7�@r/��X���@@�4%��`�����T� �N$�gљ���߭�?���D�F�Dh��Hɉ/݉��5K�nq�FN�b��&d>a�=�(}�Xe��U��:��&�痥��yRT�v)R!�g!A����f1y=�s|KW��|?a8+e���-�A�rf�SC�x�����x����uMJY
^�%3��DA�b_��C���c�LW�"��Jt�w،�����Ɩ �_ń���~hW�ԟu�f�<X��}��eB�M�_���op��G���AtPN����F���)�a�����~�b���N�o��A�L����Z@\8Kf�^����Z��,F�
e3���0����{tB ���pP���:��f�4؎QP��B��!�D��~�m�n(�I�>tNt���_^Y?�9��E?Ve�+y4�[��@i����F8�W&6�����J�gLct���o�G�@>�f�����gص�"������W�<���e��I��:��'3�ȽS����n=�1����M��PcO�ʅ�fT.�R������붵u�7���] ���@0��zZ�NbCY�zj&�����r�?t��߰�B�` :T�������ic>�c���򱽽��tםj�J�LC�%��5�v���⩰��Mh���ʣ���3RŚx[m�o]�2�y�Lz���|�y���'��e���i�(g
�HlG��x0���M�-�	{�s����א=�o�Ӟ����f;�fO
�Y)L�_�m���g�W����B�ӟ"�����bs�'�؊"cLĢO�r˹_�^�}E^���3XX�D�6� F�փ�^ɂ:sI����h�}r�}�<�ؿ������)/V���ʷ�ޒ��JД���@��pF"7S?Ey����δ��wڣG����4�|�|"����\n�n\�/��V�.�4���Eս�/D�����^+���Bxs�=e�-��J	c��������V����5$c�V�S_���M<�j ��	����
��]Q��ӯ�k���RV�+��U��q�ͺ�#ߠD���b�|e��໣���!P?w����9Ɉ/@�Kk������2ʭd{�(,
�� i	��y�WGz��bB}C�-�E��Pu�f&U�P֡~J��3H8Y��PnY��u�%���qrY��2	œ�d��C�C�\�)RM�����`�
Z����QO��B�r�I��l5d��[)�v�=�,0K����Q�1��!�� ���#�^��"wy�h�5��9�ݓA?�K�p��h�(6���L�䈀'�:L�e/ L��N�!�b�0�
�U�C���Ow#�+w(K6�`.Ĉ_4��I�L˄�Ip8�pq�Q�ʈ��j	������/"G����Hf�u���i��&?��t�B��v���̊���Pnyc{O
'G��,�^*�x�B1g�e�����pK��K��q� ?��&�ʊ,�e��}^�q�ݺ}�]�v�{<Ś����x��카�!^�>�"ڴ���@@f��H�Mw�g��=� �q�&ᐃ�NŤ��
pH'��@
��tu���3�Ά�h_����2�bN�@�k�I�]�X�FA:0�E��Q�Q0���!{�#�E�?�]��Q{l�JQ�s���`�5�A������g��}���ǣ.g��["�$���W�T>��ȇ~u��sW��iW/ox��û4>/�D�x���������W�I�}�Xjk����5)���J<ǋ.>���BD{Q��H�Q���b�*&m�Z�L�U�;��j��O���v�ri���/�i�7������~�~��Rn?lw?�)����2ɟ����B5�/@;��)��T{�.�|�.�|�:�g�O�����K�G��t3=� ./��78��R?'���<�TTHm��붶,eLaWU�.��k��_h?���7?��ݽˋ[�g��h2�I(���>��ԗ\_�Uwf0�Ȗ� hH�o������v��m��G/\?���P���R�����Q�"%���y+f��۪S��՞l�K�b��,�bA�-��&~96)��%>�p�}؃GO������>{C��/P�h�o^W�Tޤ�x�
���ӭ�f6Ƀ�xaA��1aiI�G�g5V�~}�99ѧY����8i��ծ^��6����;���T_�,K ^f��:H=�9�(|#�(���3Rli;l�bk�Ç���m���2m^*۸�,w�OΞe�3F\�h�` �*�ͨ)O����MX��;P�	,�b��q��k̥M�C/P����qDeB~����������b/�\V��ye�<���$N��FHʆ�=}*��C(��]faʅ�#��[�Τ�8C^$w�0����%S�y�)��?�I�r��Z/
0Ϋ��2�������H"#�l�4ٺ�3�6*D�er�<<(3d3�c�2�����Na�L�b�nf@n�34��D�3c8��h��U�*W)E�(��3�ē�!�M�Ӵ�(���~�D����n]�c'B�	�RGB��r�ggQN\3"{�ە��	���ƒ��k���;�s&|F�Ѯ�n�x@�k��=�.i�~\+^�\qϯ���{��e�b�
;m�=�~���+���Wn�WF��YI�r������B�2<��.�g�}��2Ȟ�5�UxO�E(���w>,���������*�f�Nۨ<(^E ��
	�xrO�GL�d��E-ڃP&�������ڊ����f��+>���%p^~cŀ=���)�b�ӄ��<	��s.t<��ߖT�74�޼~�]�~�
8���7���E�����W�����.��.�5� �8X-���({��7�s�U(�`ǎ�{���H�4��e)����m_~�a���[��W��[��z�|e]��/�AA�M#M�T������r����E��Q'0�^>,�@�Qo�c���_����E�N��Ԣ����[��3M|d�.{EW����j�����ŧw���mt�]���BT&ʕG�d�u:Y°�~̯8PF0w�z��͒�)7;��=�lO=o/��GéLW���4���8!�s�Q��/�,�Š�r�|S�l��-B�[��4*��(-��7��{��/�<q')U�<�'X��9�W4h��geN��.���I�r�o:�a���xL�dZ�-/�����db�\�-�rXn/�I���2}}t(�\EcE>S �	�!���%΄_���c(U�}���^2�J ���Ia�{,6��9����!Y� /t��4B�$`x"��t�<��0�Sa)k9���%�u�#�����1Q��W���\eC]�Rk����=y�_��Ɠ2O�d�p��
��G����D)�a��=��a��ೂ�X~�4�>�̴�)�>��?���O?��eO�D�Y�W]V62:����1���h���^�Y�&���3���S��/[��'��3�Lr �o��{Q3�7E��`�Jn>2������;fWrw"
��0��
l�O^�
���M�C����͏F4��7�Λd�-_��}��H紿�����6�^�(�� �*/Aш{�⫂��Rn��������f �>0ن�~a]����q3(�BǷ��XQ��ee(f�t^"����7!���y�q�2!�E�?:QyQgx����Z��!����C����?g�+Il�+L�J2�j_v�_�8�^��U1њ�� �Z|֥ �������mMl>z���qߑW��.�W�̞VV�Qj;KJН#@���g���W�⃕Qf��M�p/�j��q�����|����~����w���VMD��g��("?>�纲j�=�(2��h�*���3���,��@��0�0�"������؍Ke���h�V����Ud�����{�~�o�~���G������(����GRp��/گ~���������=kR�����$�^�><�}�F�ut@�h���i/_����u{�l�=��ۗ/w�#�g)�*���eO�����O�T�T�)�[��)`U!���s�D��N���HC�~������	�=��yʠ`�%�- �ڊ��e�&�[������[ �8�lb�X&n vh�R���!���w�=��c`�Y�bx~������-IYt:���0
�c�����x�i�����	��"6��:l{|�W�������Q~����DJw��HFw�@�?�D��?]�x2_��%�&r��R�}������G�W�Z!��R¸�2��x���f2V�u_h������<�B r*T�U��@���7L���'����ɝ��S�ʧ��. r��4���q�d�p�r��y�VnO���c�;қ�>�kvKH�1����C��>�Y$j���:@��>�Yd?�i��v���n
�$꾠��s�1bR�߄���� ��v��FNVnWQncE���Y��.�h���qv/2��ǟ+�m6�j #�:��ʇ����@�V�e�{�y	��r����Н�x��k��͏�QxR�9�8a�N��_��~��#�(3�!���z{m�����)+q�������ma(㊗J#@�r,���P^t֌J*/&o(�|ME���op��FVR�?�ˏb����ƙ�fDwɯ��GW��!�
H���V����hK�0h�5�O>� ��+j~t����_�_��gRr?mw���*y��%ej�=O�a��W�D~B��^8�kQOŋ���e��YA�V2���#�dm��P�cp�}�L������������}�����y<&�_� +��}�A��O?m_
?���W�/�D��-]"h�a.�=�l���(�Dʭ��3)�U��?iO�Hy���`Vy��)!7oq��E?e�r{HYQ.���������
0��ut!(�M�
�� ;�/>q�ӧ�}��"F�:�uMu�c����tf3cI��'B�)�`�	�a�O~��U�n����tNO`[+���i���'��D�/3�&I:�x�x)��|��`A����) �xrH��rb���W=�2��v���8���h'�$,��_ծ+3e&���^�:/������i�ں�R~�)�5�%���n�p�؟�b��G�c��\h�g�r8;f�Y�1��}��vҚ�$0�b����+��#�r+tއ��Z�kt|��@l/��Z�1hh�E+��%Z&NؠMgǊ�
�)�da�$Z�_�Q@������ B�%V���@эFGc[^^��-g��mz����?�|��Ppy4C���g���I�䗎Vt��g,�.D��2�i������d�=/�]�z�]�v�]�tY�-�-���N������w��#����}��F��DQ�|d^ڃ��|�Y����5�>��A�3�r&�Xv�ȼ8%}"��;�N��bu�G��<����O)��U5�B����)-�r�˅������~�٫D�.��H� ]�"��w^�$>e�Ңt߸y�}�ŧ�W��E���~�-�[f��1Oϟ��}i����8F�OD�ຼa��	�oO�\-�j��x�<,F8�C����[e��ǧO��W_=��-��7��|�X��)'\|���|�	�ǒ�%OX�$��^�c[��F��>	'py��Pn�GM0xq�ۯ�~����OM��&糓9����>)��<����(��ʣ��Pi�\-ۓ �L�%	w�C�e�6����=z�T�I�C�i�k�9N����~��3��3Ny /�t�m�)\ ɾ��/۩g(��!GM���g�y������ŋvt�Ɂ�09���P��=�@?^�VnM�$�	\�/0�&��g �×��?Ow���A�\�a�I]aQ�q&5�uڠꮑ�g`�4f����j�;Y>�/%�	H��s��گI�W��p���m�S������8	��|�|A+���U~�Ð�}�2o���ݼ%����u9������1i���T ��*@n����oBQ��(:e���4�� �hp�-ؕ;`�f�F	O@��<��|�pLs��w,����s�,�(�sF�P��x"_�V��H_o���)^r`�P#���-;%37�;��=8u��Ki!?>�xYJ��W���[���#>��A��`������"GA!����sK���U�X���UN�r+�Q�FI��XV�<���}��2����[�k�fǯ����3q�q�-jaMF��/	!����H=�H������^{����U�mx/Cd�e�2=�N%1G���,���	����*�sN���J'᳿�o�l�a�DxGv�(�Ep��{��Wx����o۽o��m&a�/�){�c{�.p�Ui���Ӂ8o��T�ha`�S~�Z��!����ʨ��}�~�����x_
ڦ��8�%�seo\��>��V������-�E��D���	�N�����~�yP<���ck�&A�����v�ޣ�����M>C.o���N/�K��Ԯ]_R"�����hV�H�},��9X����E��j��/�H	�=�o�sj{ܩˬ0Ƒ`�4�;�I��qD�� �x���#�2t"��`Ǩ��'����������M�=�u�t�l�@����N B�e�ٽ7�G�Y��8=�Z�<� N7�/�(ߏ�%Sh1�x�S�s�� m=�_�9Q���LJ�?��w����nN���k��(y�V�'Ap�:�-m�~���c�]SSV�� ;�n�vaЍ۠+��)d���r;��&d������`���W!HU����:��?2Q��c���/��Xn�PrH�t}Z�a*3�s;�C%<��� J���t�C\h���	=C�ْ�<�����TJ��B�GgcE�{���x�RX�Q)]^ �1'@xϭF�H� �����|�
x<�qz�g��J��ں���5)�Ȕ�b�+z|�~w��򣔣,J�����q��ۄ!�1p�V,�HX� �1rR��|ƫ�;>N����2_�A��~���}����5D�uo�-{����x�ʱz��%���MA�_wz��=~�Ӟ<���(2V�{h�<���=acշ�:N?˅|2��h���[;R�������ݮ^���Y�C;�o4!�m���w�_������I��e&�(B�a[��	����9��t��ԏ�Ύ�xӇ ���c<�>][������:}F����G)���/ߴ?��q��@���V��Q"o^���޽��޹*e�Wo��?%Wi:���.��W�KV�G����x����<kϟs�?+zJWe��|l�#���C|� K0��?h�Z�wH����l�Y{@�u�>�I�P io>���V���w7_��_;#�v��-
���yD�?$e�� ϔ�,��=	�5�ܪn�+�|녟��P0���J�J4c���2�X��4X�g��������I��	D��3���{p͗�$V���}i�2����U�2�\6'6H���f�_��68IFrv��x���ӕ7I g�Z�ȘJ�w�'x~�G�ps�a��]�{����^��E�D��X��=Ȥ?_i�q�>�9V�d��%�_(�-�H������ *�z����L,�"L�
�'�ۼw
6&0�S��7��gH~I'��9�YK��M'V)ن�j3g?�geK�z���A��E�GZ�pg@~��'P��D���)t�K�D�(~�j�:u�0�A��ӫ�E��	���x�|�h�
B�G|��;�q�>�� ����@t�6F�{�5�d��<P�8��/�I���-�tŎ(�5����"�@�g�u�(gLd"��/�q��/+L������갵�/e`��|��=���omʵ�мd�"i�c�rO#�٘���=ْ��nݼ!���.\��7�x�'��-*{�M�Zc2��$E}�V ��	hyD�'7T�E6��PU�2_Y��+n�|��wڭ���#_�	2{�d�}�����߳�^{�tS��_�;�#���e&/���k^�n 	�E0��2)t��N
�s����s�V5);/�,�>��Dc�}������~���Ӥ�|������RЮn�;�/��"�}�{�sE�v<g���|������l���*ʑP�>����/U�7��o��V�q�,�\��r��x)#��h�" �x�泷��?�D���T)\h�(����)*�@���I��,)���&����rX�;{^��$�uM�}�`e*|x������/`��XP��M��B�哯�5���.����,w9L#�,D���P�{���X���bK�s����r[}A��{���qh�3@����:|tL��}�+�G�)����e�5>���B�����vV�X�7�4�a�9�a��`����60�eH���.��Uv�d#���6\e���x=� �R����K��J��A,�&�]9�C�����i���Jy�#�hT�P��yfQt��t��	��Yi�
Q)+dқx���F�i�B����1���*2�t-Vx�j}c�Ge]����ؓ��~���czmeS��3�J/0x�,t�o�`�V��J*̲���=ӭU`+\�{�^�Pnh�~K}�`F�n��e���ٲR'\+v��P�߈���	�a�-�)�H�<�2;*ʟy�������x��ۼq�>��}Nz8y��%��q�;|�]��0�	)��j�@�-C��9�VnY��rKg����}�m����RNxL�ͣR�%{֜�OB������NN���ÞaJz��Y�'[��|�b��û����m�$C�1.���t��,�$�r�xH�LP��99�J��m��m��������V���؞�t�����/?n���ۧ��i7�_�~iV��lm�o����ߴ���>|�\�8�x]��Yϕ|ڤ��m
<f0N��N��Qv�b�{��83m��FJ� ��v��(�`*^C�k2�Tz+*�7��×�������R�zR�Z�P��.��)A(�ܹ� L�v������3����r>�xV!�I4'^�Cy<s�}�K���{�\�@�R'Ji�Ut���e�tY�N�-5����� � ��ȖS/|�E1��H�ʍr�2-T_�T���>{�RJ��b" x�ԄsRj9��[dZL�X�p��5p��?�$�Wy�Gyhj'��w���ho!�����z�đ�j�񲤳�^O���KH��r"<maj�s�M@%�w�����a|��E2D���K�����U����*gN�,'�՘7�8Q`&�����m�{bs�p�> �h���<P/������{�����-_�T(����"C�����z��.�n�L^��a��ˢx� ��s����.��r��f�x�v�)��L��5�F�pwB�R���}�["�=���E'D��O����$p�_���-�qPx
�V�ZI���7��IM�g:���C̼O�h�����n=�;��+���4f̴����<O)&<R����g�Z�n+��N��/1�6��Q�]�;�s�@ݏ�
4�� ?�^�.s�N�S��H

ʖ�dtӔ��ViU�U�f�) ̈�E���thf���Ѡ�1XC���W��|wL(��p��ӟ���4�y̰�I��g`��E���4@ш�2>�`�6��C�zr'��8��f2ǀ �8�x�3�^J��!>�ˋ4�n^o7�]� J�L�o��)/�lIG�䑎/VF�\�]ך���ǈ���9�a��cŖ�ƞ�"����nܸ��l?���v��e)E��Hq���	�Ǜ�Rj��o�e��-M^ڲ�)�b�ΒF�|ġ�r+��B��v�Yn����x"d�t`�OHҼh�Uh�tnE�(�礘��ŭ���k)����/<��h�k*ӛ�/{��}����V��;*zwG��0�d�����h�y�OVpY��3�[;;m��L(iJ�#��//�q|})+�o�2AB1p���(��d�,��rGV���	�)<H����HeU���Te�˂�Սh����i�~���T�Rh,�N�� �@�*�'�3�X9���ϒ���&,�Tv��%/�0�w��-��z���'�$��F\_q��DY �@XE�<��?����,�h�W;�yO?'��D�AU�@��hC�bb)�c��SA������O����Pa�X�-Μ��*�򤾓S6���I]�;,�*o���%��-����AO>���	\J���.f��&�b[�"�d���_.�S0�"��� d+A�`w�1�pd�0��u�Tb2��/#�1�a*�_H;y1vfͷ���͂���M�#-'b��U:�~ràsE��18/-Q�(�ѨSA�ʭ*�*T�1?���lxRp�1$J�b����T����'y
吼������+�h4SÙ {� ���������?B�od�0<p�����2�,;9��� ����q�`�:GZ�ys"_N��Yqʆ�+GЀ���A�,.��◹4���C�C�=Ӝ
l���ݞa�G��x�\b�r|~���������h�#)O�.��l[$�H&��r�'+�]����S_��1�UOL�xG�y��8����K�O�k{C
Ѫc�����n����7��U����>O�>���H_\�����j�XS����zlV=��A俣y U!���1&���á��~�=��R�z���I����?x��8_���T߮]��n߼�'\���ؼX�S���kHc6�ю"�� ?�y�r��I��RQ7P�v�����N�ٍ�Qڪ��������޸q�OX(p?hW��yb�/����k@�.���uP|Y���B�G�,''��ѿ�<�#�C���ܲg��(��׾ޞf�k�}@�]���9<G!� �|�-M.ħ�9q�^,����r�/".�2;E�`���rҊ~=�v���K��<���$�P��)Ϟd�Ǭ�2�Y䌟��랞��w��=�nf �o�p�!�mW�E�ݦ���___s�e��I8,`��]ń	z�x���0b^0o�UW�P�h�!+��5�<�L"�N�{]D�i����hFzoO�O��`X�H�BБ����0�N;��vaL2�¡q
	����;�P��L��8�\�QJؚ��i�'���3��C���$��(���yO��N���13F�� ��r�.�|�rJ��������G�AN!+��ė��\~���	R�s�4b�䳍q�������R��Hx�8��l�1]�k��nί����u!��2��/ެP�_.�j�Tx��Qd��ZWpy�?:Հ�/�� �O�[�Am��,����V	��D�d$yb��N�x��K�<y<Vz�G��o��_��%a�r��c3��Rn_�:Pگ���������E)B�k�$���ޡOm�����o����mϞ�]��`��f:Fj:��2��U�(���*�n�R;��f�+��N}Sa2�a/_P>O��Oڳg�l�����p�_�� ��ä�8� Ю�W�7�\��3�z��@z�e��A�郶����Ƕ������ϕ^��n\��Y+�@��b��?�[f�ze���)W��gxyl����Ypr��EU��*)��%��G$SIN� � �0�\�"��{��)�>�,'���K��(se}u�Âr���g��"�7��9mL�%Fx(Ӿpc�����1�\',�?�e�u�D����n-�"8�����:�%&��`m��cY>��Yҗ5��r{N����[$�lr�5��T(�D8�D���@��@T�Az��ER�s�I�7�gph��Y��d ?\�
��*0�LƝ��� �����_ ���c�
ddy1(�W5�T$����9��/������o��Nt 
!�4b:ʃ��\:�#��T�;4�\f�����e*��������0�83_�If�:��GE��  O���2AІ�j2��Ml�9���rb�9� Y�\�eg��Q�'�-��e�Ns�=�|����y/ᦴ���a$�e�wVly�/h��#AŚ�������8r�G�0���l��N=�s:*Y�d�.�\vN�XYe{����ob�-gn�dP�������G(NO_������^$Y�bQW]�'m�:��̡�H(@���i�"�b��>��z�]��֮^Y��̈́�rv0���9h��C�}؞?��edƄ�l���|�s�m�Kd.C�d�-�=��L�y�OH�E�����ު�2ynE���`TF�>i/���^f&~�ϴKV��[W�r�嫗�*��[�bem� (���R��0Z��&u�GӼ񿹵eŠ�=����k�9�K�[9�~&Vn{[2?��E0�nU��W<R_�3J4/n5Oު_������*��[�,/����A��N�d�᱗À�/��c��.O7��P�8���Wo��j\����h+s����dpP��F��^vX��*d~8�ġ��O<����I{�f��/,(�N �;O���S����tTWT����R���p�]�����d��K���ܒ?Nȱ�A�(øw���؅�B��R'���.7���.���v3�"A���c8O��h��A<�k9�N�PJ��	n򍋰9��G���1Q�WJ�̅Pq��,8�o�m}e�Ȁ�U	�R9�HPR�3����a��A1ae���w��4��nK����0���n�N0��GdCG�R��;=��7}N!�?+�1c%,���q�L�xip���o�X�eS:�� �$E�N�_���B��b��ōp��������H(�KI@�T�޹�+�$QlW�9wU�2�j����/��p�:���jE͉�G��4Ԡ0��1B�I{���+���Gl��
� ����^���/Vw�
��Pn�)�d:<��� #X7����d��^l;:���C���X�r��.֤ts�����kg�O�n�{��x�/ZQ>��	�:�q˪�B�Rn,[ڹT]�?C�w�9 8�n8�}�L2�2*�l�g�Vi����*���yEY��۞>yў>~�[Q�>�_�u�j����v����[6~iN�x!����O�S�h{��Ͷ��`F2���Ɖ�/_h6��"k���J�?e/�ʬ ����]��H=S���?�d�>f��VVp��_<E;��0�	�*(�S��C�Cq�!�[eۄʒvB��S�N�Wyc}Óz+).CQq���n��3��{�d��"���QF�B܄�^Ġ�?�$=��r:��ζ�}ϓ�d�qY�d��>�H,�䔆��^���<�;���X@���BY�ܲ�O�H��O���Km}�䤲ȱ@lyl���4Q� ?�LNue�<]6I�r3��>D;*,�����v�IۘN@�1���w���`��٨��M��9���2vK�/L�-�@��
����[��vڽ@��ՃD7�9�?C\Z��k��]@v��S}r���Hƫ�����
_uJ������t�t�^=Q�%�'����+����� �;��B*8|E�e6&oyY��c15��<�/I����q]vi(��y��P��~Q�.��3���[�(��t���(7
Xl ����@�{�S">	�x��Vtl١ D!<q�9�"[�l{�V|���x�^<߲R����>��]�K��y�3i��+��[��8t�<ze�d஁�_>B�%��҉�<Эm�㞗�XQ�?��	Ꮛt
�z�Gھ�����;'%pT���dv���{��\�b����d�牟>�m�l��?���>ەUVL�Y���H����KȌzJ=�
25H	;�0�Ņ|M@d�z'L3���CiB_��U�r�~0;�$3�Ĳ�i���4$���q2/��u00N��>F��U�|��n����z��6�R�)�c�B�sН3Ob��jۑd{���	����c�IR�~�l�@)D����oq������'f$�]3Z
-�a��2�e�;���>*��0�c�3�]�o���W=p���1ỳ�:����^�L�� ������1��Vɛ�p��h*S�eچ�ѭ6�����'��G�}�>�p�_��>Π�m������-�|��rW�͗|\D��}�a�9���>2!�]k̋��U�l�t��� 2��ޣ͓Y��V=V�����pȏ���3����(��q�m���O��fʄ�p��F�f�aQ�~/�|�d6�&�ȸQ�+o����ĸO�#��2b��
@�O�B�;��y�'ƳbbF�[��3]�}8�Y7g:a����#m�8�sp��;�~;� �{�i��F���F��M��
:��]bK���Sa�MBT��R��xV,F!���?w�_i�f�� N��K0�`�vq�x2@#l�0V�xȿ�@r#�� �ᬮ+�ޡ���B8vM$\##>�qo�p��!���Bq��gyeYx�|�s��?�K� ��1��s���L7r��#,v�@�B.�d#�8�eܣ����x��(f|���@����(��Rn7U�mw���YV9U�ީ�V���>-� �N��u~��踐]��h�A��C����<�]�Ģ�eG��N���4��钀�2"'�5^��My����'���/��<�C&������v�ۧRp��j2�.����	W�9g~�����h��d)�܂?۩w5q��.�D��M�g�Ҏ��a�u�F>�y��0�&��&)j��\S�6�Բ7��g~��\	�d���8J���߸��zU@]�aৃ����l��v��q�	VM�P�9��$�e5�=�����ϴ�W���o�*�J;�3�y�+����6�	_� ;��!�PF�e�
�_*S�fD]�vV��9���q$c�=&��H�$0{��Ō<â�*����&��"���鉷)M�r�����v� ��5o]q!EP$�I��m��r�pN��$T0�ug7�t����8nڎR�%�hO2C�Q����f�L�d ^�=2�;wr��R��`�<��o�>3�Ar�G�iU��c+O����J����5-Xpϊ/�:d$a�-�!��,� %@ڿm�h��x�y�4�\':�~�1���׼���R��v��(�2�X�� �Ls�����1�x���Z1��=��|@��#�ca:S(�	E9�h��ւw���:.���@�����L*3A��@�Q�lG�rrZ̞*�e/���IF~�E�[��"�*��Ȁ��*���N�\�e���{�ų����XGKPXQYSN����X-
p.�l1S*W!�1�	b$�H2.�n �nŻ�*3��}ļ�{���Id�D1���X.�H���&�a�(�6��al#@ѫ�ya��bˋ)<�f ��'��<�j8�����?�x�a0��	�~8�Vy�Uax���Y���ȟG��)������|۝m>��-+�dU���e���PQ�d@��������<��t-��Zq�4�IZ��=�Y��r��e����X]c��:�m��|�G�ʋ��hQn��E9�����?�� �ѱ� �K&�R���[/��2I�r�R�v�r;/��Ns����=k�~��{���>�<�� ��(�^�����u&�#� �'��~�(�Έ$ߜ.��x�nY��Qj����L�p4P��{��A�x)��4�� ��
�CW���
^a��G@���A�Z���BD)���r��e��^��{�H�j�����M�-�ҟ��J�ɡ�C��$��U_*+�vlgy��e_M�^��*+^��ӯ8u��[��ǵ%1�a,`����$�AȔ��h��M?�1���/�,���q/Tp���[����{~��ʛ��o4����8��q��0#�UD	Q���4�4�	�ʽ�w��`���/��Lɏ��B&+��K�]�7��ݒL�Y�iھ'� ���n�Vp)�Y�_mC���<E*������yK����pK�"�W��c�2�3י4�b|�r�M4m�=����q�w��T��!�9���ɣ�L?ö1��?}�����jVuiI�uEy_VX>a_O �1��0��{�OrK�!Y`��ry��JF�_O[��0�(����}� Y��V��e��|a)x4�J�����_�t��B���N�@/08�[����g��r���$��4�#���Tn-�L"0�	&C�vn�����G����"�/Î��fr��L��i_a�1AѼZ��N.ܒ�(��r�+:.�*�̫ L
'(!3��@� c`�
@tV(vw���a��e�*�?9t�^pɴS����Y������Da.���F��Q��Yzp��d%`��f)��!*�L�*�[fA;`�_�e&@����A0��č$�9)�|!F�����Ex�*i?�ӏ���֒�����_z)�hkQ�ܯ��H�DY�*iA
H=C1d�ho�/�{���X��O�z�)�МN&x(�TL
�yG�A������ǯ����� +��;�������:����i+�I�ŝ�qb6X*�h[�A�uLZ���R|�G�I���<���ܸ������M�E$���'=����ł�L��4;��0 � ��(�BO�s�x���@�x�?���۴]�9�3&����\�3Ya�h��K��}�¾z���(�INKx��#��Y��Ky.,��`NM�uą�aT:n;N��.d�\)7!
�xI��v���%����?��@�^��ɞ�z���8�l�:-R̼�v��u��!2r�y(�
%A�?�E�-�Ll�ǽx����0�$����e�IV�X�S"�*8+��ҡ3r<�Y.�x�=ԩ���.��*CʑG�"���K�rq��K�[9@�ٱ�L%[���8�}�ӘQB¨��E^�(� ʋ����.\f�U�_4g`p�H˰(N�����c�	�?	�L��Zʁ�X�L�\��BKP���{bR�_摺_d�J�&�q��cu�{�F&!Â�OjW�t�^0ݙd�)��aލ����/ӕMwݏ�9�)��t�����|ȿ��2�P� �_� 7�\��~�(���;�hX8�����xg��%W���;=�R�`"B�L��&Y�6^$����IҦ���YVC�~H]q�Az��(tM��9Ie�/���g`A���=���L8񿂠�k���3i��	J�K+����\��S9DbjT�I=;Bw���RD̺,�F��)b����9N$��IX�D�FU�c�/&�
�;+��P<�4���{�n�������}]Ŧ����R�$������([����ʞ?��i`�E���
Ԥ��y�{:2��c++��Q��-�/�H��X_o�Wb[�ط7_���ړǼܶm��j�2��~� 咦�e�C�Q���	�և��節3��bݞ䱧�Ȗ��M)��2�快z'�W�xu�UJ�O���]Tr�O�s����$VHx#�	
�]@���d/���S
�|Sv$ӥv��߶�̽!cw�u����k�[hPn$ױR�Y 𶃬�� ''����:~Q�CUT��F�k̤[09f��)rD9�� ��])�l����T�}�/�+b&I]��Gzu}o��J�5�2E�8�I&$KY�3����O4��hB��2W��Tq�qQz���� ����9B���Q�%j�����wLBW��ĉAGRp��5/@PJS4�A�F1�q+z�U�-�ӸXfbɆ�����dƺa�?���O�
��:!+8Y�e^�eTUL�0�1tF�"��o�8�oS�=.z� W�]���o6!�RTR��p��_	����Q�dY�x�/�+�A�8���%X�S_C���S�?`�F	�@TЃ�CJ��Uc(d�iT��<���r��e�]�6�łw��ǀ
��dB����t�v��'�v3G�����rk�b����sv�T�c�8b&T�). �#L�NN�26*�q"A��n��B�2	ʁF�r"�Έ�,@�܄��qH&���+@uL'9�#����#�V��j����'�c�@q�����
2�x����G�� _tf(F[ۇRn9�e�|�����d��I����(��Ҏ!�F��M�j�ʄ��X�={��P�yI��3y�$C��WR�X}V���9+�j箧Rh��'DpY$g��0��Ѯ6���w$F��Ǿ��m�� ϟ=�$���#�lR"9�x�]�(��B*�5���uq?[g�0!6G�_�<��{�k��G�����Y�_^��x���R�ǀ��ty�Ӝ`��Xq/q|#gL�?V�%S�q_�}�(⑯���,V�|o�j����2g� ��x� ����o���D�{��1F��XaOJ� �3��QE��|ќ�"F�w��. �!�8��u����z̤�~A��3+�>���X_�;H�X(i�HðY� m�����_�1̈���0�1�Ir����-��1�����`�Hvv����V��Q<."���z&H�p!����8��]%F�B��W�l��gz�)b�R����>�?"���1��EgSH�q0��%%�N_��
_7���&(�Ly��Y��C a��S������J��u���}V|���`Ŗ��f:�S�x*�8c̯��x�=Ӏ���:(�lK��`)��ԠR�����i��J�Nc�eRȦ��1F�	�L� �Ro���c�Ƌ6�h���Q x�&��%��%��Lc�+����z���<��9�(�`�6<g����܇s�W�-��"�m�/C�^I%Ϫ[!��Z���lGʡ�W�
w 5)�ô*e쵕�uι��b������J�Rǖ�C�*�}����Nj���D�}��~	��P�2��ط�������3)n�"��[U[���!>Qn�C4��Q�^��8X�'���P��?��oJSϼ��b�7��q�S��3C$gG�o:���{��:��|S&�^=��>����D�u�ͶK�&�c�!y�R����,�7x�8����t�M,��� #���ͮ����xD_-4����e4�u���dz����iE�ĺO�tD��vL�r��~�N��)�#��:��0��snĉxy?�}xJ�Z(ݯh��cA�d�v���
pv����,��&ۢd�܌�v����(a}�J-:��v��G�4 a,Q��\XǤ^�<p[���ps�I=*��YqF=c��ʗ�f�]ދ�'|�S(�6����������#~Tv+�޼�:Π@t*=�����h���%�ќ�i��0(i���\W4ΐo�x�4�^�&܈c�4l��4p �(�Wi�~"K�7�n3�����$�XF�{���d��[�0c��7�!�4�j��H��|���'=XdO���m)�/}�.{8Q�|����7Y�h@��f��<9L�r�x���m|
�ܹW~���F�����ﶟ�����_�����~�~��_�_�����gw}�,oث�Wmƃa�(��r?	���G�
.#7r�A?���/�rˑR �؆�\���UR�CC�D�� �p�`���^��o&���2��*i��a�؋Π��aV�f������`{��rG~�������[`��8�*�[��ͤ�͈���6�7�y�ܳO['8�sB���\��B��b��O4���!x��Q��w�rz'��$��@^�_�"�F��'��\�C^���� h���9�G���E�VA�צ���n����-��X:�{�̉g���i+M�����%��a�3"��~@٪������=q�I�/A r����!�`f��9���}����"s����T�d�4��
�L�pŮ�� ��X�D�r���6��r+p��rP~ěƥPq��
���� �f��Tq����I#%
D�{Ä��4ɯe�lY�B��p@ҏt������9�J�sك�X��L]J+&�y'�����̙6�x;t��A���W�c�%+x��v���v�҅vNJ�`/;G�=�b��x�����g�]ς���Y2q

��1J+��T���}����|Tb����{��Q[;�ݸ~�}���7?������������������������������/�������oۗ_~�3e�H�)ɇ{mgW���7Lx�ۼ-��wQ�S������m��H�w?��H�v3�e[¤dĪ��?˰������f��`��@ؠ2�'�v�f�yJ�v��y�"3&M�aL�R�T"��c8�s�H���|��f9Fj��U\oM���֊�? �](�a�t���9�cE��<��:k$N�����qw8 �#�i�y�t�pJR'y�C�u�o��Nk��aj�b�0���Q�O�&O�&�)��Z�r�BC���,�xx:8�-������I�1��y�%A���`�1�'��3�@�H�x��0���%E`�� �K�	*Txea�8�� ��$� +�GԈ_����.�O��7
�Bʙ�(���.U�D�����G'�+ l�L� ���!��Q%�L'Ҋ �id8�ʂ�{<'z�7RnbO+w(`�I�	9,���F622+;7�O��C�Y>;���A�~�H�<�Z9�Q�=��T�X��=�C�i�ffɘ���WC�V���[ŝO�9/���f�q�Q0���ݡ�'��#.u�?x	ҁPw��{Gyw0�c$��I���<�?��kˡ�(�F�%���]+���|����i�u&o�?���Og��ra��h���W�����7�rp�ƥ��۟�����~�����_�����_�T���w�����o>~&��������>��x���3J�pw_�-GII�>QbAYOpގ��]��G���
�������
[T�NX�M�H*<��C}�� ^3�̄��JVtQ�?9BHv<�4\�j[�R��=�3I�[�%����m(�y��0N�Z�5��if�J���C�����g�?x
L+Y�/6�����Tq�<�������'e��������?�
�o�]�
"7O<�1w��UP��0�jO���5``N�rݕ�--��>�X�
%�8�GЙ&A�Y�:Ly�8Aw�m�ar���i�FV�5e�t�
��aA����rtL�p��aK7[qI��28�#,�
S�N.�잺%�'������*�+�ٶCD�ٿ���S�Y��l�@#«�1��H�0$ .A��1�f�/�� �e��F�i>�}D�� ޸�`��|�BE�.g�G�n��
J�u����QB}0��|�ӁO�/�������H������˴��(�hFȠ'{�c��n��)���X�3c1y]�9�����pK(��2]�1���J3�	]�i��
�A9�d����ޖ�Pc��x�k<r���,=�#�',W�Lu-�i��%�aZ)��,�D>��ǵ��y_3|�g�e1:� >I 8"��s#�]�h��:[a)2��&��k���7Otp�>�xA�-<G�R~���Ao����ȟW#����]���i�Rn�GHN�"� �d�4�_J;�Ll���VTc�6��3N/^<��ܾ�>���7?������/�Q�������ն�*�\��/�m�/.��>���ݯ�����ߴ��?����_��ݾu������z(���kVc�k1��=0{��>��B����L�Ũ��5�|�=��S{��Z��J���O�t����!},�#��g��x(�~�3�s8����pT���&J'��E	�b�oڏ$��R"�
�2�@(�Lh{��+�.�Q�d5R1/B�D9+>�h�#���J��We3�o^�c�r��E ����k����Q6Qv�2�����A.�mǇ��7&Ğ�y?�O<�	d��U~I����˾&�J���+xIS��6�3�����0�Ë�^�#ot���G����ŝ(�P��<���S�J�yS��<��z��[��(�d"�N�_�UQG�|i��tN��	���1q8_8���tȴS�j���xj�~!f�L����f�a�5��L�0��
����2�!�&p&��@�Ic��d��,���C�ϻ��Gz��&_F:�d��X��V0���1���=�
�]n�ωX�#ȥ���A2�n�f5��]���i���|�P�H|�3X=P��e�`��l����%�8T����/�g��t{r�)��A��Q���%��q�Ü_v*3�e�V�A�	����#J���O�� �].�K����%�~�!�+'��{�<&9M�J����@,C�4��e|��W�8
�UŊA]����S�0�,Y�S���D��i� +��q�E5�Ȋ-{m߼�t�W��\�re�}�����>j?��n���[�΍��ڥ�vau��נ�,+"����/���?��~�Ň��i�ٗ�������*M\8a�P�5K30�P�G���Pr�A�,V��I��u�*L^%c����6�Vr�z�3"Ս�]_d�}Xd��.���y0. �w�+dr�K@�
jH�cW��S��S�����l��N�ᄀ�O�z?�>�|��H���b,
Y�Y� �����,��8���)�~��C���3����z�~;y(ɍ<�G�s_㮝����o�$]��9 �1o'ފ�@d��}��/P`�D�5��ɼG �qWnu. =%!��������F������=⚛���D�q'Yp�8�ʛwķiD�K<�)�k2I���٠GE���`Ib� Ү+�V��X�i� �ҵ5X7��5׉�

�a�sZS�� �D���f<R��<2�be�J������b���q�Up;�#d�0t)�c}Ŵ}�{�6?��6����y��]q~ \ N3ù'O�����O��$#�U(��B����q�-_�qjJMUQ�\<I`�3�����W��a�@"�PPp�d����]j7�]n_|�q��O�Gw��kRvy�!cY4���jB:X�^��{��J���+��n�O?��nݸ���e�����00u2T�"|��g�B
��ฉ��q���-�����L]�A����(:<�gf��fbe��?�7�C,��	c�Pd�\��؂�O��M}7Oj%�m28���i�/<�8����i�7�<2�ۂ�k�X�2O˅�`�2L���8�ΤdbC�S:R����!jv��f
�p����v��d��+�)�q�W�:���#�9*����0NH�P��PU�Z t��%�'��� �9
o���?6��{�%���*���5x'6�G�����$0%��8�+�@��ӈ�H��_7�=��'���ߙ�?���7��9�Y(z��Y�Y~\�B���2/{�f�s���-�\ G��7��Ы:3��}8Q��cq?��}Aq����˪m����ƞ�U?���cB������w)��]Z	��<?���C��� �vȹ����\�&�������7ڇwn�k���GTj5+��g�׽�YQ Vq�]^m7�_^n�/mxOq�T����!²F7�Qr�9O��/	�O&a���i@0��9�N����m(s�t�i(Kz� J��`� �bAd����ERaFۓ�C����6ټ��ir���Vĕv�����	"l�?D(G�!,s>��mAw.�ee���1���µ��k�1�	A�o�c���u2U?����W����l� B�0'���Ĵ�`��MaFL�nY�X8�~�x�d�s�ߙ���m?�B�����"Ƭ�NK�]�/W{ɉ�Lq�����U���@��qfE�}T^5���6���Nc"�C�Q2��
�0��'��_�~�]@�H�T�g��*i�2wDg��qr�`&��;��@A� ��R�e�݁p.7߇U�l�����I���Ut�vsy�Y�> ��J@q�-�t�B���>�酟��{���2�5���%�Ӕ	"�<�!�FB�kq�s��W�"�<�w��̆R��̑M�[��2ժx���ڮ]�hW/����KV`��7���C�Y�d��9ݣಂ�"����R�9z�������#��(i+���>��� ���)�ʶ1���/����ֻ���E��O�>
L�d�ׁ 3H�H{�%� ��!@����WG	�c�D���0V���l^,���?WJ��c��H����er�~r	��+�����60c`F�D ��w�I,K\��d��^�c����aw��lA3Ծ���M��@1{�d�/�X����E�i"���L9kX���L���op:B��Lu���3�3�P\���X5�sS�L�FE+<2�2mcr?��I��K�a��&XH�$X�r?N�\��C������F(�C�`��Y�Jw��'`��{"̄�z�N��
�}#�����+xC�EPq�q�:�'AK"o�/�q��;����!���zo`�OzZV��3�ocj�@?O���?�eq�:឴w�s��aF�aq^Pt��U��GUC���S�,���(�1|�H��\��"�&Z&�֟\�R�>е�����J�XG	R����IK����j�Q~,<��9a�8/�3Z^^{���r��NP�2#�cXBJ�����ڴ�dP�R�!�Ta�./�t*?ҡ����-��y�^�F na��6��f�O�7�1�5P��M!�1�S�E!^"��+?C���t�����������J?me)�񿌷�iG��c&X&�΃�[!J��9�7r?�>��/��e�Q���=u!�C�ӗg���n�	���?��s�7�܅�34����F7��ٞa��Cp�f���%����\��̈�0�7��a+��'�_s?�	P^6#��=x�fO��1��F�u�X�� ��b{�/��A���2�	Ȅ�@ݻ���$`�
74�J}��� ��8�����p` �7t��a����[a�	�sA��<�T�	g�ʳ}����+�7�t�KF�;E:� ��s<�{���?~�i��+�?L#Jn��b/ĪW��n��;���!��)��O���%7��tf�I�p�^���%^6:2�#N0��WPV��2&�i6�SjN!`t���P�(X�G�	�v�J'��Օ8{uI
�����O��_2�|�̼G/�	�v���Q!?�7�)�|5rЇ_%l�v��2�Ae$����@�3ԥ���%~o����EY��)� )�d/@�!"=_ą��$��D�(�1�ؼ���G�u�����.ǔ�i��-hOP�O�^�"OU�g��"��S��N!{"8���D�)���4�/��O��� ����u�c��X���-,���bBD�R��q7!��n���:���n�*�o��T�I���J�Ӭ\F��`�����p�a�g2��,�Ί�BJ!qUƲ�1�f7]L��ʜY����1�eh���c�E�Y��g�_=q3h7���_��<$�.0���7���h�`w�Lp���[%t��V�xH�nvY
�N2��,T���<d�����Q<��G��������%��B�F�5���2Y�������4e}�O  3o#�:���~�>��(�DI��
O�%����@'ԍ~kS�W8�ig���r�\'��{
�f��%*�̽p&�����r�M�~-yP]u�"(99Z�wT�zS
���*gաz���CF�&I�9�����[��o��ٕ2L�Y�!���V�i�<���E���%�8q̢ޣ��6�q�L�A���_̧��Ch㖼W|ˎU�X=$���Ц�
��Jn�ݖY�S�cE����ڵQ>�0�ynV�ʯ�!���B /�,L ��3tem�5�b7�2����I"S@��PAY:H�Q��J�9T݌2����2��$(bW+�δ+�	��� �"~�쾋:U�8o�c�')V�N.��@yq�!�[�t���ed�Vǭ�����K}@It�H~�����̢Q>�v�#�u��v�8�+tS/��D"��~�� ��WB�N�����e�6y�,F)� x�� ��1-��͢!�^�����J ����_���d�v�B��~�j�t`���OyyS���Ԗ���q>��nl/�W�g��:����
�:��*qh�R:&(wu�VFe����Xi�`!R9�3;6��0�D �'V��~(D�Ybv n��+#P3I�G���sJO��+0Ӗov��r�{\b =2h������2B�Y9��ޱ���f�}�R4�@G�}[��4�7�G����U�������u)�+r�\SF�r(���D��N��܊��ӱ�W>�th����8��_?7Qv�/d�e/�ᘁJ�f� �x�`7b^�@��a�� 9��yӟ�#
vl 52�8nV<�e��R��;�w
y��i�Z�%r��O\�˟�����$z��kLK�V��y ��8�]�2V�ɣ}���������y0����XY]�٦����{9����P�`�#H���5#	+�޳��n|8�}S��>�2�j�E@6"ϔ�gQ���?AY�;�:E�=A����9�(��+'~|��g�*]��H�9nJ�a�
���:e�����Ky�_��@N��e�0'��P�X���.\\nX����>�h��\F�i(�� S�47����q���v^�ɂ��=�%!�}I��n)�<<v�_!����Ww��݀�-���@�)����D��hgA�������O�I��(��9���Uo]�h'Kˑ��K0o��I�H���#�O�ߊ��8�����8=1�N�w��ȳΞz���:#ɗ�Q/��7��y��D����d1	�#O�cf�L�.��w���ӓ`ۣ~��hW���r!��]����"�f��D�S=V^����c��+hz�3��	jƌ�;Ң.�?hU{p>�0�6~��`�}��,~{�N��e
�G���(
��o���o`���?.b�<E��<q�>��A'g�H���0.:�,(��p:���x6l��Y��L�iGߧ��Cy�����]��xK��J;
�Lxښ��"����vUb�=&�WV{�� ���8����e�9��QD��ՐiVtkP���h_�����WHa�"�71Ҁ�CO(�)����8�2���d]�<�"N��w����h/0���#�d7�]H�` 0oG� ?i���@{V�_+O�S0x:R�!z�?��dX��G� "���Cv=.��'0q��H�W�V�{tD~B)!P|�����}��mސ	I#W�@y�Q��J��.���R�==�8]Y`�;�U��}��J��?ѓ!e1�!S|88R`cc�z���ENTJ0`||� ?"��:]@.^������@��+��F~�6�����6{�ʥvYȗ�?�ڢl(S�%Qd��@�.�yo��Ŕk����/�R��,[�[�~?R���S�ҵp����zX�v0���V'������.39�E+"�B�q�ρ#T����$輧[LtK�V�$ Ά�y�1'��i����s&��B�{*yE�� w��P��,�q��l����r�b��n��4ɡ��$�	
�h8��`U.Z��K@#��"N�3�*�D^��G�c��T�TNq`���i�>����R�����(
O=��� o�10at�_��=�������q�Q̛36�
W��􈎘F�����籘7�ա�AOT~�)�qүӛ��o�l��1�c�(΢h�p�\��ȩ��ʖ�)���Y��
��~
���u��~���R�_�⛰�+��agd��XX"���$5k�0^�k�~me0p^�=�r�j8�P9}o�O��,8f���K����x�K�d���Q��콲8�,VG�Ww��Vwz�0F�Ȑ�
 .eR�=��A+�erg{�mm�Z���z*hr�g�־إ�%�Vt��������v�qG�č#��8�GK8�n�����	�ö�������7��I^D@���|(7�H�HB�~O�Q�<A9�I���l���uL^�ݍW�(�@Ʊ��
�j{��5�U��W��o�Rl�9�y�ē�-�$U��/��h�D���Ʃȍ����"5�G�����q2o��[.6˾"�x��r#l�q��:��xYO���� �t��bAk��^ĬDx��r�0����o������`G�0���^#���i_����*�����*��Z~xG�Sս�8��!`�R7͋R��b����j���Qގ�q}	�ox���1;eס�w,X�6��X��&P�ԸO�cr�P��Ԭ��X� G�O<1�B�-E�ˌ�B]ScJ n������ȑ^�i�pƳ��G��0�pRذgVN�`vO��?��^�at?�J?��ʑ�F�Z1�@1��&岘�v����wJg\A�7��*WX�v��<8���=O���A�(GG�B	���W(d�Mg�&��f���%���{ ���{�l������ho˴P�{����gR�=f<�@�A��2+�1;(^q�2�o��A"y.�� �X� ��$:�J%[�h�������d%�S%��~�7(�lG@v���a���1��N��[�2���-��J.��%��M)��ڶ��g/6��'/۳��m�@����1��Z�Ŵ�u�4�ݽ�ms���x�mZlo:{�O���gz'���%&7�<B� ���r�pa�]�r{�ꕶz~��f���mn���\�.@Z�et
��{ĉ���vX[�S�!S�w9&� ��3{����s::���$M��p+d���3
\Z	�v
��x:8M����~���:͑�s`�_�n��a���4�At�v(��1�|2$�0r��������f�f�#)�O0��2O�G <�8Wca�g���Q䇏m�V�ƩP|�㶀��yX�_n��X<A��/z]�w�te]_D� �Q~�s�cho��Qf�Ɗޜ�[���Ȉ3D
�`i$�d�ן�e.�`�.�2�1V��"��ƍ�c��H �Pf<JO$���`�I�#Ƚ����Qx�Zcŋ������fn'j��y���U���T<3V�P�Xm�U@|c54�������nAp}�Fv�.��܆K�e唕I:��������.�����::����XtQN��P���L�r^��"��-�@��_Vk9wy�rg/\�K��b�h;���C���h��	E�����3��r�=|����{��{���^;BA=�r�,�Z�'��Gv�H�|#���=|�+|ў?�j�?(�+*g)��J���A�I2�<,�T�$%��g�A��ɁMNf�x�B�v�Z�|��d���[��9hO��lO��h�;�^���$`+|0���M%FT�G�ۛ��㎢6[O�Rv>���E���q+���x���#I���'�`��O���4!�0�v�.���,^t���yp�,p
��w�f&�����#�[�μ���'�Q�j�ȵ�H/�9,�ĺ��@��'ʞ�r�9?9bLLٛ+�+x�������Eל�[���dQ�g���.�r��1(%�y9	�Q�9;َ�ϱ�:`Y$��������PJH����c�D��l[Xa-B����d�)����(a��F�Z���ǒ lwO�����n'�Y�~8B7f�����rR8�籠�ǂl��+��X}h0P��uȚΦR�G�c�A�|�������=�gBu��9;���rp��,����@m��j-o��)%t�~aEaH���R�2/���ϸBy�� ���>ʤ��7�D����W�� V�-&+�K���u����9���kΨ���m
,��|��Ju�{�9�R �V<X�.-�/g��������W߶?~�]{��E{����%'�!3!��+�y$�}���wԞ��k��l�}��ݿ�L�n*�gQl�E��B������3�;B��[L%�r��z�����������fŒ���{k��=z��=~���܆�A9y���N�z_��m��&&K���-��H��ן��8��]� ~]�WI����p��J���nՏ�w?��]PQ����H���n���q}\�?X�u^��Й�;�� �!\����n��oZ�=�('X ��"�(���E��`�|��A����Q)so��&��Ҟ���:J��I?�+�.� K��~�<S�vA�;�uX�&��q*�3o�'yO,;&~<�T[���=�~��� �=��6����T���i��s�	�FGGS��*"	2��B�mn@��h?	��ؤ�|w�6�p�2N5���ȰB\�(�=j�}�ʭ��p�T�S��`���-i�W�)L�֎�+�_�1ZL:���2��O��
��%��	1�� ��l����	���S1��V.�@[A��i;m�|?e�ǛNRl��%����u佮(;��Rk�+��ͫ������ՋmE|��ѡ:)B(L>1�\���������� _�(�q����ް&\W���ݝ�������?|���_I����?|�^l�])�ұ���ʑ���os�U{�l�}{�E���{����7�W�Ǌ��R����psr�Qb��v(���#�oM����2�̐	['Te�ܶ�%�)O�?o{(�U�	�z�XV��y�Ht��� }H��6� ���P�H�b�|EI����41������>0¨���t8��Ć0x���RD���N���Lx�=혉��K����:i��0��Jn�sޜ��������ݼ���c�q�g�����άt~�%��v�?+��4�b�E���F�/�.��t�_�S���b d`�
��ƹ����"��)>����)7�RXn�xއ�-�����@~S���!�#|�e�q:����'7q�E�N;O�V�w(���6����w�.�4̕y|�N��$d�Q������Ou{ƿ`�N ϑi0mE
��1�W�D�_(pa���7��3NB��4r_�y����6:L�zFK8|{~NJ'�G����2�����D���
/ 
�' �j��`����n���I�8ѝ�=�M���_�VZ,7*�fY*B�2O^Uκa�g�Y�Pt�4�t2@/0hC� {nKP�=����v�v�\����Y)��ܮ�8.��QtgEyݽ`&t�"���+��i�v����x��^���Zņ����r�z�b�q�J�r�R[�XUy�����_]��(�%+&�ua,��GFޖ �si�҄>��l-x��$E������ @������z����c)���=����{�}��S)��o淿�V�m�|��=}������p��Y�Vڒ���s����r���'���[&u�	�/<hK"w��v��%�lU�?�r�����r�P��K)�[�PʸW�%`����F��8�R��W���6��>�/��>$�)�3�a����~_����+A�K����Hb�1��0���֠'�$�K�>N4�Pl�:�v�H��y�T����OH����ɉ��R�Mj>�~�1�`���p�6:8���or���'oeޓ����m�a6O�P�~"�p��H#T��?�m�������3䬼*���:��SW����h@�w�΋��:<E%#�=��h��&�c�FZQ����Ag�SP��m@�SɅY5�@yI�=f=f�#��%X���u�J�cfH�f;H#
t���:"�I�]�s�U0�(��`��:���1T ��`��?��;E�$��B�-K&2}\(�I<]6���^��
 t��'8��Xe����uɃ�N�P<��Ϙ@oL9,N>���7��'���}:�Η����2�	�7������^Bw'b��:@��cNI�ɦqJ�=��@�UX|d2��S�G�jO!ɥ��=�.��18�y���G��
;��cb�Mŭ�*o:wAG��h)9�T=\]�D�o��7e4�4!ϸ�
��(�o�g�v�]��xyjg�=�x����d����3m}�G��mueI|�>K��~�\�?1OC��\�	�jIAB�}��WK���Hx(�'�"^j;�-	׮_j�o^n.�)���~���:H�:ʊ.u;i���O��
~j���W�q����oK���Yi;;��o�������������?���o�m�����^�_�������������������?�����v����#���s�s����A:�kx�����f���f�6���k�+�2����A;~�}p�f�{�v�pa��-�<dK��k��A{�t�mn�+�W�ٓ�y�(�����.� C�ٟ!�ڮ}d���	\�mS�ȇL��o�T�l�n(�+��_���LAiȴ�gY���#�?���� �2J	<�NW���H����dȼ������3�,8�S�4���dɑ�B�S$	?���N�_���<�F9�/���-��Y�"����vG8��"�&`[2��ʶ�T���R����� XT�N��/�<N�ӑ�&����wa�!���诣��TCi	�QMր�*hd�t�׍l࿠m�P�`қ�G��\��t�p7�|G�鸱�ZY�/r��$��ٻE��"}�$|��pO70R���4yw����D"e�Hj��U��L���"Pf�N�;;cri���6���w��$"�+�H:�VcN�!hС3���xv���B�`5ԉ��]�U���� 3���pD��}����Β7�:b�
�m	0��id��L����Q!����<���G/G�-_�����s�_���s�X�0�F����A@��Xf)#"_��"�g�T �ˆ�:2nw��"���u9��p`��ç ���M�慼������K)=��Pu�����2��ȫ���%�IG��>k�H��P#M�� D�^1p��+�϶�����`�I��������vC�핫�ޤ�jB揥I���K	��JCq��en�Si�"����Κ��#�5՟�W���˃�ݷO�o�m��������������o�������i�U��?��߷������ۧ��WH�2�<J�ޔ2i���%�����@����[*�L���9j�����+�wo�;�oJ^����i���N{��Uq)����l��|MJm�h�8�e�LN}�=�W��#�;q�>+�|��3���	O
ՏV���.G%�q��F�݄/�A�CɅ�Pj���'���I�B�S�����gd�B���{���H�D	!O.�|���yT<���F����"KLV�)$��.嶀x�7j�ݟT���3�g!�E� 9iE~1#Ϡ=�����v;$�-Y��Uo ǟ��!.��W�;�3L�ꬔ(��W �������%���\��� ��p�ewҘ21�i��[��t���4�P��]�Ge9�`Y�5����F#�1g��r�[��AI�e�VA���W�%9��	�9�$x����Y���"{���}#�;�=E33x���sNc��U����ǃ$������fQ(
�Vhx�v ���� ��J��AIb(r���'�F®�)�V�=���rP�aoU����P�y�����2r˩V4�6��-�%!p	�n`5J?�|�ёQ@gF<1(+lu�,P�.{��⛭:G��'�Eq�ʳ_�b��|Wz�@	�O��H��W��48q��S�v,������a����O�,�P��t&�tky�n�#l�0!0���_L'�e''��������#F%�ո�H���xY[_,+kKejz¼��{�Ʊs�bv��Q�Ƌ��H��,~�q�d�I<�W�����&�a;:6������H��>-�^n�xS��ǧ�_��?�������m�~������v��>*GGFA���-��[P$���/Fx�Xy2f����ӧ���:�vd�}Y\��Q�������Z��X���xzzQ66w���N9>f0�e�7-U^��%n���zͮ��(���P�^�̩ɨ����:�*��Z!���|itC���5�?!M��2ǘe��0NNN�<eҗ/ćtr�;����LɁo��, z҈:��D���7t_��6�`����y��T~U��S�l{�.�[���fd�o�w�!H����/$_s��0�깋�AY���z�O�8K5���+�_�E-Fg��ʈz"t���%���"�RqO:9u�t�}dؙ���sݨ��i�f�oM���;������?�|�`�rD�l�JP(��)B�<19aE911aE���{���nI��x�н>�!�����K���UZð�� ��E�E��Wiѿ��м�����^i'sz0��W�����!��L�G+M�z�n���I�S!r�M�Z��\��"!.����{B(.Yv$�4)7d�l2�����r�m ���Nh���ƈ�[>��{��f���<��~zv�LL1��������Bm<sn{�ꖇxwxu����]���{b�uT
lb|���O�{�Wʃ�eye�L�LYN�8�"���`yP	��{hR�X�$'�'��������sS���˻���������͞�[[eg�ċ���T���'�,"coۦӒz��"�^�@e�uP���܈�Rfd�߻�R=�'wE��5���]��VF���]�q�8��_��T˦<���?9*��5C�	):�15zCxiⵌ����$�	�Y�$/x uk���w����s�������O�4���(��F���<�$~9����~"$9w�=�|�ܪ���ޅ�C�8��rs�Fd���ۼV~9�[��>�yxd��U6q��1�";��`�����,��'�lm0Q_u5�{�	=��xgW�%f\M�ߍ'0�,��W�
F���C�� �����G`7���.���W��r�'ꆅ�B�>�'�_�t*wG!��,4?+j�l��`UE�N��(s����l��c�%�U�aiAv�q�9]�{�V���ۘ�{����-#�\=O�7zͧ�PRT芾WD���CȚ��N��t�kWń�N�I��l��ZEG���=�$���P��~� 4���Ɖ�0����|n�兟��j`'-7�1���V2n�"F#Jٛ
�Ǐ�w7�6E�Y�\//o��۽��/�N&Ic?7{�.������ۈ�'��!4�K����9]�>�Id^l7�� /ί<���踜����\ɸ�)ss����{��/ː{XVVV\�-gH݄>C�G����GB�EY1��Ϋh�>�2 �
#���yg���bFa�U'愳z�VLl6)�	=� ����b�ֆ����~���<����7q���[��ny�ݨ�1Z����O�/�xX�V���4����Ƶ���F��W�������Yc��8�S��9���ſz�l"�W~��0�S6��3eF#�H:o�<Ѹ���� =I\�c^!W�������)���_Э�T���� ��4n���<Q�n^^�7�NT7NOO�&�	���S����"�%� ��A����K���w�62ː�:t������K�s��4��C�I�a�F�Ңx���x�� �
~������{���`zj�x�_��zD���1�"�#�&�N��q�R��x�8��tӟ=�`�zV�ٺD����I40x�/��ψ�o�Fm~�TǏ����01�S!�Ƶ���3��T�(� P�UT�Z����7
_�
F�9tzz���M���I)�Q���pANTˮ#��]�����x4�� -P/E^��z$ ��
�]��h�a���9Х�S�!N�M�b�����>����)�5�����#*�-�d�-�B�}u��S"<�ƞw�F#������q2=#ٙ�q;=%YbZajGJ���(W�  ��# Z>�İҸ)�g������9!E���k�+�޽����h7s�yM?1�X@���u(i�AcѕO �Qyqq�xAʖ�!wjj����˰]�˸],��k�TF0��.�/z����4����(�Y_�^�;d|�g�z�^�#�ɝ�����e�
��VbqY��V�qKډUF��)3Cqť�;y�����)s�Se}mY�����}u �e�1��a�e����>�a��-ɔE�5Q����E�H�su���	7�*�~e�M]�ʹ���̴�n�Ϟ�*?�[4r*2Gn����qL�ƧA����B�I�]A�mزhѝv%L�#�ONj'K�-��������~��k���3:���>ћ���	�-ꋯI��N��YW��������tD9z^��Þ��.ԃ����y iE{�>������qU�O���:�q�Y����J��'a���q��+)8I�����k�Ի�@�_��J��+�!]��G������N�ۜ&ΟN.����:�B��W�@�ҫ6��Aa
��s�O� +L��1���V<��B�%�J�BFZ��T��5
���M�\]c�M_!�zK��=Aًsvv�LM���s/�J�h��#n����5_�J$�M���X�S�u�����F�$���}�@EC��Г�'@-�(O�<6U=�'t�5�'4�P��a����A~��k$����d�:߫1�Q�T�����i���(��$�l�HP�H2ĕQ+��Ԑ�Q� ��:J�5�[LU�ˆF 2U�$�C�Ry�� �n�[��S�t*#�R����K�r]Y^(�z���ܨ4��˄��.~��bEd��
��Уa��^F���p9<:/+z¬`�vX�������݅25�����	(fxʗ��l�*������F$�P����Y�]-�Y�+[�����l<��Zv!�b��􉳋r�!��`ě4�{���܆����R�?/�����l3�����219iZ9��Qyu\Nʾ[d��|c��ʇx@�G�״�c �M��ƕ�	�Fi�$#efzR�=�	ϣrw.���-��~бi�`���$9 ��@��Ǡ��@|dZǘ:���E��A0�ONe���Çq��$h��*� ɩy!�ø�#��z&5�Zf=�B����p�i��l��*RqK?�E�@���~�p�A+a܎b|���f���{p|��	GD���<��#S^����Y9�ޤ���y6�?�w����# 8c�t���밉�q �e�{Gǿ>��p����q����x�@�3����)k]�%gwAKg(�γ�)Gv�~�!#c�2C"���f����!��`&�P�
�0B�k��g-�w�@�y�.�n�}N�H�W<y����t�8�zo��Fh�٪(�^�Ŧ�9z�V�#erj�{r2
@\5�I��I�&�n�`B���נ�]؆���L����<I��/�*�&����t����n�I��@C��8
�!�؀h�~�y��*�=���������E�Qf\�B--�
r��-Fi�*1�<z��� ���BcҐ���\�#/a�Ĉǭ�~vvY�����1�9�t(�e��27?Sf��xA������7�a��Ix��縻���Dٳk����hc���j��K���DY[g�t��[_�vSlA���V��nCN)@����G8�\T���Y&��xw�z��w\��˞���s�jH0���F���D�oAF�B��g!��a�YJ�G�,�8e5�u��IbŸ�~�3����M}�=���07�A���A���l�~��d]�!r���L_�z)�~_�gă����W�ʷ_?Vd�{�2��BF�����wp�m�8�C�;a(olw�^y�G�ȣҊr���2a�4Q<�U��Q�N$4r81����tY\�Q���0	����'�]����[�4�,C��TDX�¹މ���guSt�^��5�\__ʸ�_�������ى��.�w@O�wa�B��㞞�*�33�L{�;Ƣ��F-mK�>�N�.�}O�rK���F�sC�)�#��*hj�n֥$ޞ�AF����=/��P�3��:ӭ���cϺv���?2_��tN�<��x�t����ByL3}��Q&ʾ �Dt�d�*�Y�*��?�k�פ������������-�.�N95yLy��L��@b���<u��s������9��q�%>�/o���cf>���d�ԭ7]NB�Ŀ��� ��1j9�F����Dd��2)�ς|j��y�@U�J:�&�~ĝk����_��>����{
�KV�T�-���N��5�8���X��E�o����U�����(R���V�M
c��6røU|R>ą��Ba�7@�<#R�4V�����g�<).>}ݟ�p�HPa+cQ&�4 � C��A�`;�M��B�C����8��/Q(A����,��f�����9j��m)SP�q�_�Ȩ�1�`/ƹ+�����K�S�Ce1&#�Q˥�)��%�u㇀�Ñct��o:�'�%/]�T�>��Di�1��Q�9������'�ܒ�HoL�;�0W���Ĵ2>��F�ґ4����5y'X�Z�
����"ǟb���#Ut�Y^Z�(������Դ�6L����q)���-�.����H^�����{�L&#��lOԁ|+����ݲ�����[P����XY_�-�/����27�Aa�����a�aF����y�J�r&��a>���\yOVЁ�g�;zy��j���~$c��mc�i�tL\�`��t��Q�d�+e~���Y��8+���GV�?��W����_����\�	����}�?�)'�ǧ����-w��C���O�������>��z�����x�*�xn�.�gzq!z����h[p����o�]�w��d|���#���G��hQB�
�5)��Yr�P��yо}�vT<���|kC�S~t������h�-GG'����8���P�%����4��h�M@}�ubbl��,-�{k�eey�k9�5�v3��\y�Dt���V�k�Q$��]ƒ����>C�Z�rt�5��}�D��{�)�a�c�z-�8A��;��llCq:^�����oa�vu�]|�?_c��kX���d Mz����5ke}}�,/-��I��R�?_�(=��T)�����?��W�E@��	}Bg�v>FQ�#��W\��Yv�|��A��(?�M��y�4	�� |u�kӅLz��䜁 �oҨ�8�/����	��5��G\�7�q�#� ��Q��7�5m���=L����%[
v�V�x���J8��`IL�F�[��xo��qF|@O�Tcp�X(���i�W�xL:|߸�L!ۃ\�үx�_ /�8!\*�(@%�<1Xr&�V=��S��R�4~�yG�Xa��M���x����t����5.I#�X�L��#>��2L��A�K�C���5�q�w��� N��d��wE"l�-�F�t�<�a|�L������]�}�O:t�h((|�%�
{!���$�'+�5��>nBC�id:�5}���@��aA���0��0�Ԡ��+�H9����P�q�� �e�I`loe�q���&�Of+oA�����W[��/�D�d�r��m%��MM���ř��Ȣ7Pb���r4R�_*!�?я�`L���Ϟ"�6*Հ���ŵ�e��}��W���9�q���<�奙r_��ÇK��;5�i�3�܎��,��-x��)?6
�؈�F��� �e�c"��?rDj�%=�I���Kz��"��wx�����cj$f%#�K�w�~Q���)�|è�J���P�9�C�-���/Ϟo��Ϸ|����Ш.t�J*�.@^<V�՗X"a�+_6�9����`~nJ8����˙�pt|Y��υ���y�D�q;�q�p�斮Q�����50��WiU�&|	@��Ж�a�4�|��@ە�hw�gt|�}@Rg�bH�1
1h��c1�$�`F,��C7���[�;�WJ#���Q�Dj��n���u 0�NL�k��e��78Έ�������/�"��W�|�.=�u.�F�~�%)��4�隤5�����C@\�>A�@2�Q��	�����p�Sm��[y��K|�m*���!1yH���U�2ܽ��z	7�]���!�����j�'&��������VwaҘ�/g�O;rk�B��n"�p��g�@�͕�H.��:rk"-����#?�I/F�$�/GG���+L����)�5�}p+�ܜ��.�����9��~�����p�0ä(���
C�0R���������S��jzTR��2o2i�p�O"p�w�!��4 �Ղ�r��
p@ߥ{S
�i��0�Ez��Ł�M��4�	�6�P�$����b4�HG׏�s����B$���a˧�Ɉ���aR=lF�9���u+֠�B&�П1dͣ��D�r�SLEp�[�0�]�7��1nO�`�k&b�ѽ�"G�2��Ƙ<ٰm���H�`?	P�W2^�HFt2����̆��Ξ?ǲ��s,~��5ۂ��=#���c����%��w�1d!���Ź��{!�x��|��D����rT^�ڒ��]�|��x�<I�#�__(_}y�|��zY^�U9+_g�����NQ #>��	��Ǽ����=����"����߄�C�����(}O��<������C� ��Ӱ2����.��?����?|�y��8��U�ޮls������_��~����y)r�H�G�)�@ؒ@��T�Ζ����hu�ʕhz_�&ƄA��1�=���LON��]*��6�ô��*!]��.���7 ������A,1Ǣ7�3H��8/�K+a��.wy8<e����(8q�u�#i�7��@�`L�1�g�����S%8Y�:OtYɰ�R=
����R��^{܀x�o�qo��nk>�E����Q������Ё?rM���8�y�x:��I���d!"$m��3��#������1P�WZ�Q�}���k���F��,�}o�8�.G�忕��	o���x����SFӭ�^�����~h�@���:������?�y�@dC�W�Bu���nB��v�F܊���P���kE�}G��n��6�<�Vl!��cTF���>��~hé�ُ�����0?7ZY�4���H��ʑ\V�{�ҚO�0���G�8^к0����Pih�M��@��5~�� nvO�i�+����Wt|Z����k�G�T��H>i�����O!\o'� tq�;i���rgd�y�����1�t�i���p�Y�$OQ�]��\^�� ���0ri`��I-�[өF������-�#���U�6>�-�g�NP��烲H��1�1��9<:-;;ew�Н7x�������� L��F>E��
��2�rq@��#�FC^�ݼ6g�Έ��Ȓ�H0��ؕQ�����J��{||�w���d�/��W����wPXZ�Q]�����X$�L'MP�ѐF���OD�36n�~���A�<�(ӠT�7/)m���7�~07?W�=X/�|�u��w�(ߏ���j���S9�ِxvY������2l�����/g������)yH���8� �U)_F�e�2��-�y1�4[��?����P�<>�c�1�
�s�k"���|4�j����<��&#��/�7�)`'rzd��@�0����ڠ��~9�{����R� ;n;�!�qѳ�S�qK�c�<b�Ö�Q��B.�##����]�X	��%�C�1G���rǸ��º��{�2d���Db�{�a��F��H�QvZ�:��R�=a�n}�y���g�FE��y�]o��)8��|��{��v��	��=��/��EG|�[��*/�n$t�����qۅ&��
w�;ЭM���,��'��K����C�@f0+��E؏��T�)�
�x>'�&�a��N�xV��ٸ=<:�E7TT
Bq�K���@o�m��!�*3�~�|������Z�0YB�Zy���4*NG�+�v39�rWj5�����F����QcŖ!J�0�1"�3�I�ʿ��Pac�8�_��K��~���-����������ˉ`|r�jm5��c[lW�B�|�S.�y ؓ1�qy��x�}����J�Jp!exa>%$���ƌ��	�&2�k��ҩR�]���]�O��5h&,�(#S�e|bJ�#2��d����#���@�K;3;�K,|�X����F�ę����dRy��\.Ut쁞�G��Ϥ���l�v�T޼�*/_n��owe�S��&F ���ɓ���wO����������zg��h���<?7��?��h�
T��~Vc~t��q]ƙc|�|�����������,,/��0h��P�P#�wxV�=S����_��Cy����SJ[e���	Ň�$^��T��>�^F����B٨�� �1�1Ƈ,��3��2-�a��L ��p�����:,;֧���@VyɄI�	��w=����I"t �:޸U����g,Қ��-K��e~n���EB]E�b���sͧ�Irj�>�1?��}��N��Y�Ρ��]���5��A�I`�no�}ш|�w{;��^�>(N�|7(������g]wZ��б$���Y�E�V�oc�pL����8�mI����Ԯ��KW\{�ߍ�w��gpvu�4x�R�b�t�="Z�A]�����Su�ϥ���rt��%ξz���*�F�r;�TXCFR�j\�KB��C�l���Wv'$����������:q�=�мHѬ?� �g�9�>W��N��[Lc��/@��^���4���=J�8�˽kFX|���h��ݤ%��3����@�p�&c� ���H����׉�>����J#�\9>��&�j ķ�y��P
��e������%X��4L�b�(U�jXQ.�#y�`�l�2��6���L�+��J�Ҏs��i :�J�n�q��Z�Ư*k�j�u�#���3b�&��YkS2Θڢ���z6����~�x�Q:b��rQCyS���[N��M��]@f�'��Ҭ�P��A�s
ʔ�*f����G�4�\��İ�؛��U�Cx�>�W2�9	l[�f�����lV	A��2j�����Iy�`U�U7���C1���?2@?~�t  Ȁ���m?��+�Q����L�N����ɗ��_=,���xdSJ�d���{���go˳g��ƛw>�bat~L�-�Y�1�����.V�8��	C���R��/��rR�{OŴ �=;_��r�o���T/�T>�i�����{ɿ��4�D#hO�'N�J�����ʲ��9Ձ1� Y�
_2��_��1z!��N�ݸ{Ӿ���
�P�X��qK�p�P`
P䔬0���x���X4��mN]B'e�dz�Y�l���N�_ܷ@j]�;te�3�NGHF�1>��/8���� tN��<���Ⱥ���3ى= ��~�y6��;@�#���J7�������%�O�����B�����S}�q�r��15���yt6�9���|���aӍ�Ѥ8�x��O��W
�k�ʼ�H˲��Vw���iQ��/CD;����C)�J���16��У��}7L�F��hf�"�D�V8C�P��>����"{�����4m�w�2y�ah�7��ň�C�X��h% ���B�{����X�8DY�-!�Abpa���W�(B�_�nMjx#��3��BUmį���JW�oݪq+��׬�ߓ��J�Y���G�V��h�Qx2�A�:�Qi�/��K"P8��(%��0�a4\��P�(<�oۚKZt�(1f����,{�N��|�W<�(��yl�?O��q�)yS�>�S�Z.~��z�?6�~��eee�;0��Ѻ�+�2"i�ĸqP ��M�U���F-��FY��?�)��:� *+�!c���}��W�>}%��O�b)����B��e�����+��OߔG�����rq&���p��c>"��>,�����~��u���`F�E�Zt����V�rnq��߿_�?���Iu��tF�1z��z��PF�vy��Q�m�ee����L���Q<�m��k�#���ǡ�1W����.d1���,//ȸE�ՑR9#K'�2�9Xbg����s�����u�G�+_*�Ӡ5�)��׿�[��}����+�1�cvf�,-,���%�ܢ�I
��(�t�ݓ+Љ�r,�$�@�C*}�<�����_j�B<vp���g���!�8����l)(C6ڃ��<��Q���>��[ �;rc��n�v����^�~d����w��̠si/�H<=?c�#�:`ݘ2D�Q�v�]�=!I�C�V� 4��0�p����5oj?@�3�����fG���n[r}`��{v���q9��x��n����<+Ըr�<��_̑��~�����#t�M���� ����8A���3n�X�-�A��F
�SI�^����l1���4"�|R�ݑFƟyu��s�O�$/;�4d:�;����֢��������]��UK�0Ղ+L�����d���V#�����j��M*$;������\+f�6��{S$�0�\� CY�l��&�S8|r�FlI"��U���Q l��mn<�h�'��xe���y�Ĉ��d@��kĀ�|�)�q�3d1J3=�
�q5��W�{�3BFj�/C���A�#�,Ǣ�g�:,�:88)�LM��Ĳ35B�9&c
�vum���/��	F�����K�h��\���D���ƅ{�Y#/\	���2n/.o������>{�Q^����QGG1�L�U^__(O�X/_~������z	�;b�����D+/I�gC��8~H��2�G
F�U�4��kR˹�yϻ�ȾʂN���Wo��?n�|[޾��dЫ�2:���,���4+N:���t�!�/l^���zĈ�d�H�'˽{�e�ފ�ic���c�쉶w��ݲ����g0��ݐ�CnB��?$���S	$r0��Z_S�\/��C��2=9��f��t��O}`����rtȞ��և�u,,;`����������i.<U�i;B��1�y�6��F����^Ա������wޥ����B�� ��t���!h���9��ƭݫߦ*�'̵f�vBy����<���o9�?��)�c����j���L�b��
����4��O�a{�rָ�#:�q��Ag������ �?�|����9Ф���7�m�D��qm^T���@�ȡ8���Ϗ�8����`�F������ �Ox
I��Jg�n���K��� a��?�W����φ 4C�<��Ϛ���W��>�w`�����(Zg�
^7�ȵ�B�	m��S�qS��3s䱋�%-�E#SPH�*^�����z1©��4|S�=o�;yZ�'���KF���0��ħ��$VK{�V�
1��T�VPl�Ι��ǉP�Jg����0��vɇ�BR �.���@6lP72��d����R�݅NT�RF��NN����mTC��{R�e�/�%�4��$E��%�ع��^���IT���4�꼨g�^*1<!�7�9�����'���	ہqJ�A�i���^dԎ���i�Ud���$��S�ҭ�w �n����1��J��������jp�ۨ���+���d����&2�|vn�ܿ�\>\+��]:��M<��F��iS��z@ܬԧ!�{mL�v"�|����3���l#4�8r�[[m�?��E�����ֻ!,�	�yrz�,.��2���dT�X��y�S��L� �2�ة'Ď롨���Ql��B�.�R&1~��|6w]Ua�u���Ӌ���v�ӟ_�����߿,���བྷlN����eȨ���<�L�$	"����%_&�����G���Ge#�7�갴8[�<y(9�o�<B�5�R}�v��-;�\Y�B/1g�N<B&��W���<}v�/: �����3
N'��=x�����ܩ�؍ ���ѵ�������/'�i^\��2�t��T���a���<��1���l��#=>���@؈��
=Lo2M��iO���P�3Mv)���H��Щ:ct��s�O >�	=��a迱L@�^9I�T�S�&�c��{P.$�w%`�8�\~�c�����Z6]_��,�t��֍�.��9n�.�-�0� ޶�d�#uv�"'rW4�jܲ������ԩ���vR_���cCY���F���ku��E�}W�>1�G���m�hD�\oLo�o7&�bE�����n�����E��:*J���|�}�ŕ�H�DwAUk�:l�d2�A�4VF�w#wܾ�i�,����4�YPm�6�L�%H�~�z��{�i�,¸M���oi�eǻ���W!��������]��£�� o�	��6�yI&kڑ�CP�`����b��A]�칫ʇOϚ����L]  ��q�)��}W�p��7�V�T�<;�7a �h5~�М�5vwm�y!��
aI��g�����<=r+c'JY��B�k�5�"�`D%��Ѡ|����d�8���Q�1rŨ���V�����R8Jv~��� w�Ϋ�M��]��9��(M.ȱ��n��Q�mD��M��(��Ėw�WV}����|��`���[*��sel����}�O$[N#�I�=tۋsOa��t�D7�2�od������A���W��~�Q�7ov%��n�gC�73&w�,-/xA�
EGJ��:KG��`B>t�������^�E�X��0τ��z�=���/.�����A��<(�^���S~�qS��K������g>�d�2: と�d0�M|�A[e��]P c�U�h[�8�a�)dԖ�5�����C6�_qظ��w{��]�ȸ=�a˗"}�h'�A�0�`���D�{�
o�N}�aԶ��?��sFe���WFk��N-�[�h)u���22�|ϵ�7��.�e��"K��Ǩ-�h��&K`;��.=zv<*E刿�O�Ãѿ4x���5�čH�X�� 1t~��ȴO��H8hS���c��Y9=�sn�.FnI�$3��˺��SG�*�d�������W����]�k�R�a�Y"���³}3r�� ���I�_J��E�`@�ѤC��g�W����Z��)x�g������s�E^���H�MHo<��X�'�a���C��/k��Ʒ�]��CA)��t�����4֛JU��On���̯�#}Oc��=����8�����C�QI=�K !��DӦ��.A��u/۟/��hM��o@��6�D���~+�c�ݽ}��CO��*�ϡc�-=Rb��p���^���(�pnhM�J:�R!�0��ֹGC���㔅 U
�rŰeq��ܜ��i�������k�CAM�������?��1J��!�2t1J�.��b����,�	 @꿑�Y��%sFύח2"ȓ=7`���\z���yGX��!�T�q�Y���dܞ��
�6!�{qa�S ?^��&OO��$Jy�q�� �sy�v>�L��������^/�"���'��G~^<S�������?�?��Yy�Ig��H��1��Q�*��Yy (��+JSV&���lU�^#]�2�"(�2f����#�!�F�^>���O?���/��o/���_���s��������,��qe�iZ<��Ɣw��2t�Ta�`�zT�#�*���f�y��p�ڒ:��-�{��˲:?̻�������wV^�ޒ��N#w���"�L��[(�[P���I�;��,�oȲ�\ёe���mlS5ˢ'��С����m�,����ؘd���W�ߑ�mp�~+���:�NЖI�/>L��BI�2�&vK ?��Ў��x��$��w����ޛ6��/�o����U���~�e�`�����J#���_�<�L9�^�
���V�;��n��ï�_��b Y�e��0�S������`��ޣ�J���fdXGK�J���6����0⃇5��o�ʻ����K\M��ߍs�Cx�ڢ���g�����1(�a�B�����eŬdF�+}����� �w����!n ����m+�ĮԢ��4�**�2�ۢ�*Mr$(�	ss�OM��ړ���ۂ��?*#��OD������=�l��?��c,���p�8���0���k�	���s�o`�C���\]�x��p�e��R턲%Z1�c�yqq�.�i av@�X~:t�T���+��"e��/
qgB���G�V��15��"��|nV�	��h�z,�Ca��"mN:�p遾l�P�N�?�ic܎�ˋ����=o�9Q��r���N����<=��
&�����6���%]��q���:&6ro�j��(2��]t�Y�q$.��s,#j/^2=��yy�jGt���W�I�^i�H]!W�	PQ�}�� ���妲"�i�P�H�cDnȝO��y�Q~��E��_���������E��_�gO7��ƾ�/�1r4��{lE�L�bGU7�]�5v��!��Ayh������ue2r�Xܻ�R<X��2� �a�6;$��>.o��躧|a��rA�4ց�Crk�II"����K�$<��J��j�1�81nكua~V��yϹ��Q�����}�	+��٢�R��I�ō�e�1MIםp��v	PnO����`�r���O���bn��,��⋏z��q��C�R�iZ����q��5{!B��؅������''�:� t{��i	�k:��eHC3�q�z�iN�:"�+nv�E��>w\��c�P�+�0T�qxmA�݈.�Dw�QSCZ�;:�9�t��y�آ����H7����#C���U���y�t	�L�(k����6�J����͗|o���� �>��h�>(WJ����$�JB"��/�dc�����w0UPLG��TP��mU�ЂວFM���Wm����H�1<�������!4dH`�C����@F"s�P4��PT>-g<+r��U��TZ}���t��b��#ϥL��;���yU����b�$?��GjK(Wvy���/�+�nм����V?B
�5����D8_+:n{%?x�^��F����C�Ɩa�4�,b!���h�7
�߻tX���I���X��U<��+�a���d��Q�yq��ekk��5�)����8��������zYY[�����	�ˌ�P�h����Hb����=�-P���.���t��Ou�Ƅ~�����??/O�nxA���E����^v{��a��S�O�IvQ�8I�s1��@��F�"�	DY2��Ex �1�ã��w��1�w[;��7�^��e�>S�7^��2ʈTustJyS'EeJ��ӋK:P��DG�xY�I��L��v.+X��"�U�����/���p=T�ay����G~1���˽�r����r��f�`�U�J�{���D�$p�5&I�����C���iSX�]����wK��+I�
S67ޕ���uѓ���C'D�w��&� ���aK�����`[@���b��y�~��l��#wb����Uz\�j�{ʗ� v�5�������.cx�]��*w�֑�xA�݉����\b`f�o�2)�P�js��F:W/�ۧ�ң>�P�Pe��E:��������27��N�R���u��A�*�v���qL_�٥���}���� ��6_��x�}nQ��YqO��]�{�[v�)+�	�^wD�d��Ah#���[��2#�q�_�}�_o��$�}�A	�-4&�j�[iK�W�Ծ��:N� d/>�`���'�������E;at�� �b�s9�f�#{�ܣ�B� m^���("37�{3"�_��@��5no����v���n�ޱ���M��h���TY\���8F�U;+vh�=������D�`�C����'���h$:�uԻ%,�ϔ���±����_�A/q�4܍�_��;7v���0�bd��'޽��"=�Y;�����1�WVg˽�tf��bh�c.s�U| ߓ����M�<U�[��x-
�X�~��E���Ր�on�"����e�xY���/߿,�^m�ÃS��R\&��u�� ��Qd�}��_���z��#��Y�"ІK/����J�흌Ľ�c��^^�/7�Y�S�."^��J+��bD#4�"~R�t��&7�w@ ��W)�����ג���������)��b!��ɥy�n�s���¨���ty�*�M������uѕ:��[�7��n8O3�,����'˂:��ˋe^�]:u1]���y!��-[�;�|[��02m��:�V�V�B��y��(�r¸E?�?,���	:�1��T�^�1_R��6��An���6uFߛ�G=�ηe�rR�n�9��rp!��+X��*�DXS��#��_�K^f�=�G�&m��W��>t��w�ޑ%��;��y�$/i����K�V�QZ]_��/��\�KvD�6��v�nh��0.��/���#���[B{�qH����ǳ���_����k�����F��P8~�ڛ�_LJ-���I�Y�aD�u��0� q��E��A�?W�B�VJ�ϠnTB�N+�9��UP]M��z����UE����h�Vi�����oJ�<���&��ybT8�B�U� �G<�{|E�̕@�7bV�L����~	��J�����7:B(�?��u�t-���@�f��|T����_�5C��NH�+䣸d��)gF���ȵ#���k5��eeέ)�`�����e�)�`:�6Q�qVP �ʨg\��ɶ?�
�!�/J�)7̷�?dӾ?!c����*�#c�R�ceee�,���9��Oԑ�i%9(�&�5ճ�4��W
��q�� ��E��29�\��"���o˿����������������)��_��d�rw���<�������J��2�-�A�r�<s!�a��0�qœ��X��3z�H�<�v^2��Ձ�찻�GG��oR�d�ǚ@�_ң��_��R�`t@D`��K�˒��j��D�	˧q>�� _&�i���ڢ���aМ�r0ȅ[�ۃr�j�Y$H'��h��䈲����R7�$��Á��F�32����5�#�~����Θ������e:��=���r�`�q�^$��7X�q���A�0Խ4l�Q�̢<�'�qp��eTY2���ɅGm�2��`:n��H+���h�{ޙ�^�yɟ�f}͈*�o��?cJM̿fWvx�o9�xJ���d� �Oe�'��'�6]a�`�; _�����0���CG�թ��EQSO�$<`� w]�>���X�?�W�?zXV������"��t%ZS�n��n�F��"*��E��Я֛�o'���s���8b��{��~��|�ޓ.Wh�nɧ�z2?}28�z?T'��7�V�h�Z�y߉�Be��j(��i ��;q����r��ǵz$h ��6q�������xb\4�y遲	�N�	���5>hTcˢ���a5�uէϒ���Byd䖅
�k��0*�Sd��~WA��rb�]a��&o�/;�q��Ҫ���c0M�I��N��[�|:��A�*�:2s	��:��׋�u�6����� e��f�Jòm��ᡑ��( ���H�ŅY��NH	�qXv�O�~߅���@��%�+��~	�0��uoK��/��d>+sp�>���|ii���@X�A΢>+G�CF��P��?���뽠��Q/q����ON�m�nn�x��8��O�2��W�ac�b̬�͗�Y:�����=����t�+ZM�Fz`�}K#I���k�\ڱI��"[��H��^����ey��u�����5��< >hL�[���-���X�>FX0�"���4=�y�����߽FʘgF�1�cΰ�*u4���z���M��z~��F<d�:�΂��� �L���h�&WS�LA)�B�K邛23���e}}�ʘ{�g\:�6n��%C�ee7��9����[�+��~�7� ����R~m��j}��Ve\Qs|�YX��BH�1�+���	��]x�`�
0�[��L돫l��� Pb@���Y� ��7��	u�c��(>��CppxV�wd��`�m����S>@���Ok-o~�������t�g�㺬6 ��������y��2xB h�kPY���x�@�isՁ�{����s��t�y���>?�j(~�~��҆3%���"��Tٶnfn��K_/,/�����5��O@���S�>]���O����<���w`��B(7�z������5��|S�ŏ��<��/��ӳ_�_���$T���R����׻�/'^�|��
M�~(���3~R���}�Ž���	��Z��p�S⊴s�u��x�3e`0��a��h��A cy���C���饻��/�bΟ��,�.�IA�������͈NGp6��+,نW��B���7�eo<�Q���i�,�Q���@��w䑼���N�����6��?�1��*���H� ��oh81`���0=;3.��f�KWW�w��tҨ\�O(n�Gx�X�L�?�Q�n4k�5N �+��c�-�o�kv��]|�Sczvq^6�6��G���[X-�\���e��?�u�C���U����.��I-��'y�?�w�y
w*�#�NѰd�fh���q���b��~9a����3�c~~���Η�Vˊ�R�|qzj�r��T6�H���:+�]^�#w
��7{��~dO�<~xxZ�n씗��ʛ�]�^�"bU��<q��/��չ21%C�=oOT��yI��O����a�b 3��t=r�Ɔ'���
�22��#9ÆU�����A���!u6߫����ZȂB�#���N���gR�Q,.n���Ɂ`��6"�Q�mYٙ�ʛ#U�+���.��o��l��ޫ��):Qz�Es���Bl֏3�/���u}���e�����Ɉ�m�5���+��A,�Rb�d��\��ɡ��<S����ۢ�<WV�9�{{g�o��{�t��<��b�Y�g���P�;���P��*@��o���,D�φ���te�����ι�=��͖�e� {�*��ʟ≑�s/L<�P�,����Bg��+_m�9�ROt��F?e�#"SȔ	�1��WE�8(��␝#u�XP�A+�|�&�!�샮Z�ܣ3.0�U��+�c�Q�^�`��As�As%Z@�aP|J������̲��8�6pQ��6t!��s��0���P�(gE�n���#~C���]4	��F(�=+�]Lwc�;O
[�_����dD�g��*�y���Vծ�x=���1��2>=Q�&'�9!ZA�E���Q9�'J��-��Ѿ
���b ��<A�m�.m���(ރԩ��{���!��E~ή��&�i�-�.Hh?��L��&�{�@݃���&7��{���p����s?��d�+D_f�~���/����=6O�,.@�!n 06�L�Z�!�gN��oFd� �0���!?<tP�T7C罯᱓���c	L�7��:��¢G�g�a5�Wj����գ�!���d�z�l��!�z��QQ�e#^ܓ/g���w&"@T����ǁ|���������'Fr�*浐|�'�9�T�e��`<������xF6#g��"��$���'L������J|���⻸�,G����v��#�J7�P�w,S��&�����s���$ m^�ЖE��\7�r��04"?	�'�s��x��'��4�'��I)S�yue�q�'l!?	�u�}!H�*d��d�+?ч��UE�sV�5h�),���c�v�l`��za����(XX����Ç+j�f�+�ks�c��B�E�#���Nr�c\�S���!�aU�����GN�R�i�n�2JC��N����?��7��Ա��`rq��t���k�V�%��~j�~V^�x�>�}�T�^�1�W�Y;�b��B�*���#�h'^w~!5��X��Y���u�_�(k닞k���j� j�cۻ��㲵uP��������n21��&Ձ$�p�&;4�L��%�,�ǚ��a������W����x���i7\J���wg�y��x,�tl�?!�J` �@�����=W=[U�vÖul��8?[� ߊN��'�Q��A�a��)ʷ���b�E���*{!��k+*�k/��eM)x-r�6�]P\�PRL+b��݋��&�/�+׵�y��kKY�k�ǟ��!�9�&NKzH;y��v�`�����r�/�h\&j3O�/�2��L�)�^r�lDZ���ga��E����"��)��5�Ss�[P"� �_)@�q�YW���;���Nn&b�ڎC�c�����9HحB�9�ᐿ.���n!�����J@O"]�ý�����|S!"�����N����rL'�&��~q�!h�����[�����Kzp�c�-#C�v��?�1��*7^>��ab����DU�;y#57�R �&�o�w-�]~D��C���Q�,�r�u@���a�G���9�2i$ȧGM��y�O1��������٠j��?(p��T�m�r�8����|�'k͏��#�M����G2z�����H^�<�t'--W�"�C�Wp$�(W�{Fav�1�`C��]����ct��ln~Z1'L�{&>dI�j�*��;�d�r7���F�7(W ���D������*t.�Ȼ&��9C\|���̸�����W����<��`������9�Lcs����]~����~-�D���Z𠭓�V��ati �����!b���
P������ۡ���;�|�Y7�zt7$����j�<u'0�_k�/���ՙ��RV�	{�`���-�Q�z�x�
ʠ�(o�0����lza��#t����������Xvq�$�Oq��n�e�FK-:���LQ`+C����c�U��c��
>�sh�ť�i�+[:v�G��:�7~J�dq5Mq���W�lyR/���T�y���Ke��n⑿f@���{�,�-�Z��tMa&�n�\����� �?!���D����Brb�&��&��)�F�A�'��ut��!�8��8�J�H��>���89P.|}e�������������#����n��ۓ���_S?���Wa���s���@��ǝe�i�Pt�q2�mi���o�SЄm�Ig�/�ɖ!}t�#`2z�>�8Q��x��8�	�;�)F0�ջ`և0IpI�S��9u>��O���+$t�ɦ��x�{Or����m|���l� !ތK<�'a���}���qB���/*2�O���x5.S/|���{Dq*O*�rϜ��kw��r P*�}:(l6�\	��x��!��-t���i"gBv$`�ٸ�A>#Ü����aht��`d��t�9��yO=�wbf��~�x��֦���X��w�zz�ܴh��"�q���	ʗ��k ]�O�--���n�τ���Ed�OQ��8�i���޼yW��HaN"40��4�Z~���ŗ}:մ��4���ԅ���!'
�z����D�t1��X����?O>?��v��4������:�k\��&Er����Sņ6�0�	y#�:m�EdޏU8���8����{emu��i`����/{{��۽��v�;=`�1��-���T���È>n�Z��?��[[�O<b�&sA���k
�8���*$��||�� �����n�[xT�3����
��Ī�m|�W7�d��s�4���H]_\Z��e!��7��좜��˸%�f@ŏB�k����"yk�C_��W�	=�=��vY��LoE<��8ҝ�we���$�%�{/�2�n���P�aĊvȨ���ls��<1���g�3E���/p�^���vy��m���R�y�),�?�(�׫�N>��֭�3u��㡉'�-/�jP�����Dɹ��-h (�DԼi�9�x���.��?��@1��@$� i�� 6�-�v}�L��;w<��6s��y�H�˷�K��3yK[��;�@�Ǔ	j�9+�Y�3����i	((я�G��O�9�M%B�cH?������F��`�kܷr����+圅NR���>�z0z����nǼ��4���P�6�A"r��:y�8`�݂N�#����/�T��o|��\�2)F�/=�������^H��F�9a�͎��H��@�<��=��Y>}���i�b8s�F葑�����������=7��6F�؏sa���8!���\]���A�fP��Ĥ���wLȻ<��^HY羍�O�o�e[�7o6˳o��ޫc6q�:��'�7�~U}q_FĜ�a�5dB��� ^��|n�%jع���>tâ[�n�Mx��������&���	@d�	CN���0�x?b�!V|/]C]���乃�<�]���a��Ӂ�3{!9��H(�����C���K��N�c������ɹ:E������^��Ѻ��b�А�=�q5����Y�yD��âU׫+��^�)���2���������3�gص���Ve�2��fv�xn<G��A�5��7ѱ��)��B)H����kT�i�r�����F�r$��:�ұU�У��p�wpP�y{�d�줌����SF
���(���u�|#���3����l��)�����D��>�Z�� ���1z\	�=�E�Gg�{�ٽ��`�;�1�Ϟ�,O|*�vS2~h��_�]��<��낋F����&'��6G�)�ʭ�)[�^�I��y���R�4��3�I��'�2n�w��OO<�Y���.�[/3�]A�<Y
�82ֿ%�40��\Z��J=5**1�5�#�)�(D�w94<pgټ0?T�P|ʟɋL��-�A��Et�$cn��70?<���� ��,�b:���Y���uP��~��G:�\ȵҌt{���N2�-ς���L��h0m�zn��PR����dYYf.k���4�`wß�$�e�"LL:+�w�;�*䫀�5�����hT=D���g�i�u������j�75�� e:6fy~����C˚�T�Ǘu�b䖆�O�Ò�˲���W2p��)�޼SǎE$
�[�Z�#y�<�_��-��ƈ�P�[��G/;��K�}*�l�7�~��y�C�v�k��ӯ ����L,嫑�.��2�1[����H+���FmE�e�g7�-�蠄Q�n����e�)�+K2j���V�ɟ}?�a���ll���v��7� ǈ(�'y��`p�q�\}��/}E[X�#�������2ne^Rg�N�5 ɸeZ��ѱ�;�^a� �"����`����픥�ڿ(�@�&�:�x�Y�������	2n�fø%�b��̉���Lb<��y�Ur)�F.["��.64���9l�ו�8�@��w�Bk��>�tҩw綁^�}��G96�(_�y�˘zE`��V�݃[G�2�������-G��#���E�'"�b�>�:yq�e�?�g#�"���s��s��@�����o�D�.5?��	���g䶥2<���k���	�4����~T�4�"�� z��)�hќs���Ή�iV�/yeS_�����U�?j�yo䝄��h��;;�����LM`�GΈ�ʍ!ÜPFwb��J�J�6��"�Q�	�K����`��V��Y7��|�jpz��kc�&+\�lв������d0ʸŖbU���Xa�-FF�C��5ʶ�����85&�Y�������Wc���H�y�1w�P�f���e�|ƨ]Y���cc�N��U�Q�� q;�N��=�t?�FbC&���Hyψ�+Ƈ�0������/m�n�J>�b F��x��6[�xr�<~t�	�]_3j{�2b58�����-����_	~�t���_�4P��蕼c��_�������2N�3R+�Ve7b�c�Q�_�ۖ�����Q��oʣGe0.z�4����}��?-Ϟ��ij�_m���#Ɂ���F:�N14�yi!iNL��� �M<�.
㖺ȗ�koa�"��5���fU|tlO�n�+����/��6�Ҧ�J^�6r+&"h�bo��EH��f�����M.�Эq2�&l�
�:����;SY(��Qӫ��j�y]�m�3�G����椻��2S��/cJ�t�$�y�Hh�+:�̱e���<s�+�i9�_z����:\�/�Z��S�-��=��[�ess����{:B��X8Έ;�Y�E:A���]ʋ)	"����=����[��_�����k\~��d�&^n)֧؆�P�q!����#P{ud���}�_`^�	d��L{v���6���A�6Ҩ��tGT}�Dե)br�5�v�8+D\�Ʀ���Pd���5��/£�X@êQ>�Q�w2�|��h�q��};`RH�KS��8����A�+�y�W|��n9�\�'	��>LM�3�W+��Da-4�7��xI�-(�g�ʧ�@kL����T�HG��D��Nd,yZ�ʕ�e��G=�5>��AQy��Ay�n"�}���#yt�{��y_�#�����#8��Kg��0'�F���T��`�ܻ�,�ٮMq0:W�vl�\*���N�mN��I7������ǘJA���)c���H����z�U^�x+C��oO�ɔ�&&����Ty�p�<~|��p�0pi̙��HZ|�C�raM.�t�l�큶D�Kb]�|1������w�<E��3_+v!�)�q���-1��9 R��ҋ�i��.��h��O��C���Bϒ�!Fl1loN��
*㡲��Ⱦ��Iy������@�σ��ߓa��힌�7����6�n�FC��͖f�oЛ�]_����3�K'o�U��@����C��~x��ƥ����ԸGk95m}u�̱eä�zԩ��?�g�8�zl�8��'�z�蚷MQs��Ab�lUW�/���Ly�2S&Я���zwrzU�E+m�_��B�Fyt��u���ԃ䳢^�}�S�Qu���莓�X<�LA	��2�pq�h�G��C|���/��Ad����[
��G���9:Rd�д)�sϺ��F�q��b�����˝rvPc@�Z��yӋ��%�U�"���;��q?:~�7�h��:i�	ݤ �w[�{A����y�w��6��Vi�h�<�N��37�zj	ǽ��`ס���Z^*�6
Q<U���e�1�i��8�k�3@���^Cga�a����:ߪP�v�l�!���6��a 9�fa�h��+�f��
4����,������ɤ�0���ב�H#����iu�*0��[��Y�����`��rɀb�P.��'+��w�/��$�T�ԣ,�@	�ͣ���7�'��1��'te9�s���!?���އ�����	�Qt:S��3������)Le�ߥ�㲷�_v�w���X���*��w!��r2;���u-�{Ū�rF:��@�me�K� ���q�����U�[���c�r����N>q͖:��������ʓ/x����Bq�cO���JK�"3;���g�6���N�l���s��'��2=�������F����b�P^`��X�x�^���Ay� ��}Z�Q:=���t2?�E;^�#Zچ3�O�	�Lt8I�z�n�0��p��.tc����B偫�ٯ��r���U�u�?I�᫩l0�eԁ���%p벦ސVM�/�ЋB��޼�6�u����ш���aF�ru,��H�{�r��Vo_����?|[���romMF͔ʎ��`>{���"s|�|�v��Թ-ҝ�@��~�ߨ�Ű�q�U��S�o�	�Q~#7u�X�Ɓ:����ZY[�!��R����5��nW�㴰���B�	+�Ӵh�iR�12���)_x᱖C����| \����Fg���A�Z��rv��#ˇ�|��q(�<R��I8h.ɵ�e�cLF�gD7�_��;� y�|f'�E�S������1��e���n��k�*:�LG���矘���|t�5�n�g�ZX��1r�ч��rhQ��h�i�� �e-�Tr�W�ǈ���LZ7:��fʅ|���1Nd��kݧ^�U���  ��9��$��q���?Qp�������W�_��DA���h٩�j��hG-C��g`Dȿq��>V��mHW��GnD��"�p�����|���6���P��ɈA��oTX3)
'"��Md5^�-��n?uӫW��O�7����H�̈́s�#�?O8�����DDC�
!�ʼ����2�-�q1*��'��K�}�;S�L[B�w8n{0o2;�J�y�>iL�7de��-|����b������v�`/A�Z��^�l��m� 7�F~xE،H����[<'�^Փ���1[ϰ�H,`�:cj o�[ʗ�HE4�(\�������t�떙�}S�^"V��]#Ge{g7V�^�'���N����e$��e5�3^�#�J!".˳��=S�B�e��碉{���O/��MR�1���!�77���e�~�������~���ciaJ��R���G2��؝�a
�e�<?1b�@'��NZ�_���6t��S���j�9ä_�AW��Ðeyy��.9�@~������xo�%]��ۊ�5��e �O|!�U��b$��s Y;S?����������<zx���=2suYʑٍ����Ͷ2���a� !ˡK�@���+��3�*��+\���Ku`�}2ᚌF���B��������mG4�cy�!O�kD�<�+Q�/�ðFF��I˹��5�}H�?1h��=�h��cLY�ʗn8>W�ԻذG,��8`�N���I�� �7t���. k���HT�yOZ�o�8DY�)b��E�L����w|�����a)�ڑ#��d |�H4�0���.詳�� �Йj�U,��Q�΄���R�L:��1�ŗ�/�G�Q�pUlr�x�!F�D� �Vo�e������/�晛~ \�# ���r~@�����ȇ߇��b�����nm<=/{!��0�o�h����7�`Wż��"�x0�ǒ��!M��՝�a�"�x��ط���@Aѓ]�򟚞���������]�,��J�����?��F&Ҙ�N:�O6bd��>����+[/XP§�!)�Q/a;����2��UFBPR�C}��oPŻ���*&����*����N�ge
��.���X���'�=�̋�c�e���X�I���|�ȁT��W�hoF'y�P���w�H2��)��\s�
!㖨������@����ۮ�/�{�+ey�3���'n1��჈��.�IDP��WҴS �\?�0���*�x+5�1�$Fp߿������^�ݝc��VJ���11]���I����H�=�?1Μ��rr�2^^0��<( ��䏁�ǳld��zaD�:�D�v�K���� �w��MLy	>������X*f}��i~��L��`�a9;=��Y��/��ڰ���{��e��E��Q'���:i>fwK��1FB�Nk\�	zT�J�E�忉�� ������Ie���k���I�8;V91�bģ��֖���ta�k����My�~�]޼a�dlǇ���m�/Ҋ��b>�b�ݖy져�����#;2��C8&�rܶ��E�wL�����[���;[bDq2T,�%fy����C�f�۞�-��IެE0���^m��jt�)yxS,L���}������W6�cp�.h��+AS~���?�=!Mt"�mLG`�fFƥ��2��`M ���D��Ϙ�è�Ұ� o0n����J���4�t�����3���+����7�&���9O��� ���%f��/i�!��x��E��?D�� �]�0n9�q��Te�N��c0ăQ{�ȇ���,�>W����٭���C/��Ul*/��9��G�2b8�O|�2�CVOv��ɨ]�"�qK��ҝU/ג�H�}���!}�Ĩ��'�1��B\�l�:�M�cK3���v�;>0oxZF��Fy��[�k@R��F� ���� ;�����# �x��vJ`�-ۂ���ܙd���f�vee��9�ym�vR&|	@�H��]~�z������mv^������,���%�6f�{��]��!� �|t�F��X�o�'���wO�72p��_�Q�L?a�:|��� +E��<�c��R`�57���G�f�� KS����X���Y�� ���:��@^�h�k5�4�`}cJ�Ď�t  ��IDAT	=u�wת/���.��/�G���c��������!��d�D�p��۝m���yQ'M�"�͆�y@�y���F��	��.v!�����8S6�D����b䙯��u_u����̤�G�}|��C0񚽛�v��qlUF�1��)i��j ��t��;��[��{w����ښ:�2p�tЉ��n*�2n����Ƿ�x��#r��q�z&_4�4 B)m,?�wm��S�fgf��pFY����r|B��:�������m 2_��Q��ˬ�`���[F�gf�=�͆����-�?�f������=(?���se��E�aK��jZ<5iV�tDgH��q�U��p����L%
"�_�
�,V���b&�G��5!����yJ{�2�#l��q��|~nN�CP���#��"�,�<��T����;���3�C�2�8"#���?�'���W��Q�ɩqFc��9�)f�JF?)k���C.w4���e�B�=<�t�0-#q{�FCwvw�0��sܦ�GD���V�N��%���P�%D^{Ӯ/hD��c�Aqc�ҟ2w'�F�caȨ������n�f)�/��..Mʰ�_>�/��hN�	���j�VrA>j����wD�m8h���E��b ���*�'4���OQ�x�ÃX7.>�Nɨ�)���_����c��?W���IY�a������3(�.�Z�@�F9$v���-FWt�½^�O���w iޅ
g���!��}�M�W��O_��z4	�?h5Zv�b�)�d��^6`Y�`6��VG����W_�AaSf�� ��#��W��<{���y�]vw��=��{���mEk%9iih3�m�G��,��W�V���|�~�q�,"{�����V�F��0���������ͦH���J��?�#1W�#��{��_��H���1��2⹸����ZVW�d�;m�;���^�މ�a�a��3�Ms�����C��}Ӆ��� ��&H�vWB~��Qs2�3��.�A���XG �v�l2���o�.�jZ2_~-`����*_�ivf��Y�|�=��g�KȌ�֥�ț~�ҩ�N��c�6`�U����灣�F�iZ�"{ȻQ�n��AQ)AW�%t�*t�i%!����^~]��t���C�-�U�P�
=6V 3Z�\-V�#��J����q��R�tv����hF�� ��� ����>)�8,9ҏ��:z����*���\~�vZj�X�J�4�m�GY�G+%��Oʋ�#mb澥����A��w<A?�{�v|B|g����gǄ�w�ƃ}� ��L|g�6�g>�G��^�qpL�i���箉�(F���t�w�usS�� %@ڿ޾�)I�����r����eu��9���b;4QY�%φD�
4�	��<�U�v�{�5��[�q���иd}DrV�=]��ק��˷��6��#���M'�ѣ���=.���ߖ�����'�QO�ob�%�Q��S����߅�B /a=U���= ��G�w+|½[�z��4����X��)!x��kb�N8�YQ<p��>���Q[F�d�]���8]���a��w_�o��2�x���(�0`��O��۽���7���מ�z(�(ua]�[�A"�V�B%�8�n�nz��3�d�{>S0J8 eH�{҆"����_�\Vϵ�^�8�P�����fy%�e�$��1Rbf���Ǽ�t�BqG��A�il�٩p�u���q�fF�-s��d��ɉ�8򪬹���=P'�}�c���:��m�Y���������qx�^�kt��F���'9lc�!��8������}�am���u)����y��D���&?��ŕ�iLa���9�zA���lȨ:�ωq�_��1��#��܆;2|����Ox��Yء�T�ʰS�������g t�ւJ}�������b
̟�ߙr�_��9S�m�����y����57I�+�X� ��y
�l�e�>{D6�)yXFߕ*�y9���Y�=5A���죈�4<̈ �#�R�h� W�^�@gtlTH��­����E �>��*,���9����-���!p��m�-��(3��H7���@��狰y!����x�SD�r�g�!V޳=F�xa����Q���)[[����1:���'K��?�Q���M4�H�'B�s���2��`���������WW�dN��E��� Ǹ=���-������iL��4E6�Z��|�|�N��\�A�#.�ގ�s$��k5�����?��^^��.���W���|���ɣ������Ͽ�F�ja�T�5c��7#�$�A��w޷>*��w0Bw�7����RDϧ ��9�"~v�z>./�Uq a`���#��?���V6�g��Ir�a��UO�����B��ۯTn�+�ӕ��ӓNg��޼�Uٿ)�ӳ����ʻ�=����N�[a0%��f������s�]n@����1��G���
��2����8Pdqq�#�L�XW�1�̞_04N�z����$17��O�� ��7����/��Y��Skҽ�Ɓ�8���ڄ1��G�3�K�l�2E�z�Q����M���a��Z�w�[�e�t7 S��~0�[t\M>k�t8�!]!�_(��S�2 �|���S6	�ƭ�q@��Ύ�V�@�Z2>�a�p�!_Q��������p��b?�9�D3M�y��֥�����ݬ��K�G2��vL��C�FM�@:�����w t#���y ����ȨDa2�_�h!㑯�<�����w���s �	l�"��'D�Z���t[t�:hZ���	�K�zʌ�1`(Z��+��t-���K5�tN��a�ː<n!^&�ܐ��7=W��DD���<#>��FdTBϼ�q	��e��+�D�#�H�ɟ��8�̎z�pb2S8n~�Q �-���2��M{�Y�?�w0e��:�
��*F]������z���%�ţ&F��씕2\�Тe
�m@+w`�z�Vyi�1���y�M�d	��S:�WcZ� �X�e(��c�/�����ѢpB�"���u4�6��P����p04EJ|A��[���@�§��(s�w|\�?��##<�ӣ6���K����H����N�߫1}����Uj�!]<�ǖH���4���2F��rL�`�P�1}�f�<�<�Q^o��cՍ+šz ��ˣ���/��y\���aYY^,7�V�r����(���*���J}��K����z(w��f��%� �w�s���7�.9��~����;�װ���|Wͼ���}�,i�89�L��^��%j'2X����xy�pŻ]0b�՗,
\���| ��ޝ��/ʏOߕ�O�t�]��Ine�^�Q	Y%�l�Ħ�6jI�0�lz�.�_PrL'��ӆ	GCq����_מ���_~��<y�@��l��t�4��I'��mg��4ꠍ.l&�t)ͤO�4m�:ӡs@����-(�,�8���V��3ݟ�S}�6b�,�.3B��d�.����p�\���H/p��C�d�� �*QߙHa�+A�)hg��z�Q���Q
��1�9u����6O��o�'lav����u�����<�S@��H�� ��xH��0�6I � ��~'P��O�VY{۸���23)}K��|�I���3���]Ҥ�=��nUVy�T��+8;<W��J��	���Y�!s䕯l��*$��DSE|��v�7����^!��[浹�n}i��zj@0�Í_�G�7a�_rs�j�u~;�?7����ikQV�ڸ��ddIB%t&;z����U�d�)���7�K"p���4\��I����ˊ�Ľ:�_�H��p2����U������Y	��{U��r��5s�8��������TY^f�m��-|���J**��1�A�?�Y�����J*|uAų� �׏�\�f��'/��F�kE7@�lLϺJu��G�S�Y�@�+er���,�e���&8�H�z�\��B��"1{ܻ��ţ��f�$�;�k��H\�E�!.���f�^�ED1��c�3b��6_��͕�9>���#�vO0ʽ�p�1�%M���b+��	�=t'
�̝{��<&od�\^��#�����y�F�DÐd�#��j�WWg��*۰���j8m<�Ty���Hc��0R��Gn!݉��p%����m*;g�f��;j ǤyzvY�ll���.��ey�r�#6(}�vw�$;�+s���ߕ���O�o�*�+˖QV]3ZN�@�y�[ӣ�^�eގV���S~�)#`�'l-W7z eآ;�0v͈Q�N��J<3��o�|�Mr#�z��
[��^(���<o1����*���A��dlݚ�~&��:q�͞�WWƱ��<T��}y�h�����m�/���7�|Q��V
{���T�:4�/�)���7ʟ��Y�=g_i}��	�W>�_12�T����k��}��g�7E�"l�7�u�	Y�Q}Q����E�Ǥ�%[��7$y_R��������(����
���bwvOd��Jw�9���F��3��:�L���e�lĨ5}xB�p���y@���hbN3���9$/���H�8�L�Kw��0�Y��(���+���w'2�D��Zl��Kp(�-&���Ħ�~�d$�������\�p>�g*Ȱ�5;;^?Z+_|q_:i�u�'tnNN\�d�z�Wŧ��b�E��yo��st���ٕy��>��SQ�M��1��=�uC^�RS�����ڸ����[��K������{�Ӷ�  u �3��A.��*���F����h��	�M襊�f��~m>�g�U�<�-=�n�݃ȧ�P٥ma=�2�)�su둓�D���`���t�$�G�m�j���{ΒA�z�W�;�}ȳ��z!�IG𚠮��{����ơ�d��7ėq6����q|���HT�[�7���x�) �n&��!�D}Mp�q���^M_}�G>�ʅ�X3)>���&sTO�μ"���4�y��SR��!�7�_�|�,z�m�k�><�7����{B?�[�/0/�!����a�p����7>�3���ȒVP�O{�' ���H���X�!�D?�H����¤����h��ŷ6�B��(�膇M�GTC���hFuhc4qee�ܻ�PV����<;ZP��HD�Z1`���4u1����1(��sUG0n�G'E�X9�q@û�qP67cz�!Fs�U>q��������	ҌO��{+��~J�1�2u huD���)�h�d��'J0�2�3�9�<����k/"bӧ�ߖg/Xǩk��OCnf'ʓG+2:(k�.�(�%���gW��&��� �؅�[���k#膉�E����'�3
����BvA��?uX�\��o�N	I��*�}����@1$f���@o�ԡ�IE
#��'Ǳ�2FWVfe����8�V���e��a��`��>-/_�?�Y��8�a[=;��qW�c��Wxc��|���j���)����UP�)���0�:��8���=�]����<\��~�+�I�]�����qy����Q�0����ΒC��0j�ϴ��vG]������S���(�rFn�e�NM2 2UVE/'���V'����nm�=�{*���䓽Fi�j�F��L|���to0���}rO���/[aܲ�[���-_��i�j�1�Lۻ������<�jz]r-+\㱡1��cu��=���.�Z|�F-�zR�9�6�K�,�f���̴��	u~���7�L��	_k�f�Hy#8�~�e2v-7�w�H$��j���w7��
�}�'*�[�F����"T�<��s��g��S~�Qu!��ů�G}U�N���K_��r�l�4�̂������� ��_'�@�?5�O��5��]n�0��Ǥ�b��B,�IF���Y�#2n�'M�!?B��Tc1��-S|�9���!�����=aPV�n�R��h�d���y-7Ec�]���t>�]x%1sA���@�MJ���`_`��	�c*�����B0�!
�P:�\�3n+��ŏA�e��E���Fe�-�N�m��yC�_�e�C������k�ϐOj�##�ڐ�Ym������G�>簎�M����jT홷Sz�F��{�`0G���!u�&�@�񓵲�6W�ԁ�ԫ�s0�)�STy��c�A�C% �MO�O���AU���^�)H(P*��1��G�b�|�U~��u���7�����#Ye�ovzX��Q5�|Ƭ� +RFLا�!���/�o�w0�^W�5��u2o¬/�?�!8h��T��e�����]������E��AW]���W���emm�<|��<y�X�㲾���Y�Y���ۻ(O��?���ۗ.gF9��N�G@'ԑe���.1IJ����?m�8�g��oŞ�!��FZ�h�)E���enn���___)�3�V�Fu�}x��°�x�{���c�2���L_����)�˯)3�I�B�EF�٧s�I.�)Ð�z�>�A��ڒ�ȅdW������up�o��`Gt���9=@7t�-�y!��p�׮sB�MF�h��mz�7������Y�!^�"�˚֤0����`F7Y&H#���v���}>��`<��7�u�z��ڪX��@��%e�(��̌��ϙG<*�hoE;�*��ڇad(��>b%E8ѢI1�]��6��R3 ��#�֏Yרl�M����ߤa��^��㚷g�BR��������ŏA&�IH �� #�$������O����ip+������Ӝ���a@���h���|�4+Zѓ6n'�v��ۘ�@zT&��V��xV����J�U0��0p���y�/��
#��j�G�Qħ}Fn�/�Ӿ�8�Jc ��|��,��%y�#�F�׸}�]U,= �Kx��Ɨ�M��gyX��a�����q\v�ʊ�uF�gf�<J���zy�`]eĶ`ʻ~Q4�(��b���������+6<a�I&dl�x[�w����0��|5��N����:_�?X��%���[�ݰ]���X1���ō0�3&�'OJ��(�Q�]�+���U�F���mn��/6��?��!�Q�ʐ��=�dćQ6䇆��^�FT�e7c������3� σ����^�N�Aއ�B���O��N����C?����l���^���d|r�휖d�/��������?T�vc�����򗿼�뭭]��d��c�i�)�j<=��u��Ԅ�G�w鷃��kE��_��%=G5Cߜ���1�~R��e�{?h�ėٽ���V��|��i�F��#-�S��H��Y�+�f��~]wtkz�C���o�;��[����M��\^^���
�<� ��Zȼ�#,qr$�u����g}���MŻ ��T�ǋ�5���:�v��@���`��̳kΌ�7�N��1e�]���+�}���(�����"��U�'?t�
�4���o���3�!Nt;�#�1��ilǶ�!L�l�q+�Eq��c�E�̍����Q�/ �����\!�� ���x7�N9����(�3���z3(��c�?��}���p����C��H3t���4���>F� �dVW�zap�W�6�e��_�2Fv��u�)���Or�����2^@��@U�����A�a�B��yD!yNF�1��A~���ڰ��7� �;B8��@���a9:������@� /�Sϝ�����fd%&���DK��H���~{/����� ^�O�*�_/yq����ӽ��_��w������3>���dy�`�+�Y��U���^��m`�>3實�>�	ι�ɍ���#n�+̂���Co����g���\��Ccfv���-�/�xP>\����j�9Q�'�|T�R�,NQí	���h�r1B�mK�|���|*�_^3���s���:ESjԆ�({%��?�*��U���Vy�q 9�*g���x/C��w��!�rDVp=������ݸ�Q���@>���Q�:����ti� ��4�������QB�1��I��/�K�����céY���]������ߕ?���:.O��ޕ�S��`cZ�Q�H]o��5�A�l�ϐQ�r=�Ց��v�P�ٽ8?��K/lz�����@���R�\H�X��v㨼x�S^<�T��uǷ5J�p1㍤Y�����QMaO]�k���`2}@�N|����ə�9���w����:M'bԝ��3:W�����u�t�qY�A%�u4\C�k��P���#�j;�>�-�^����%�v��2��;�f5A�1dkÝm�&�W����W%���W�EXq��ԛwa�\N ����Ѩ���O!�O����Wo%73��t@<p�����6�-@9�#꜎Ieq�:ͷ+
TW�'�T-;��p2�t�H΍�<�O�V��g� ��^��D^̳��7r�OZ����[�����7':xܝT���^qY��L��D�-�{��2H8r�Xna�"C�$�|��V�Z@e��G385F�S%U��O�FmUNv��a����Z(�;"�W�!��?�bbt�����?R�嵌�8����絘S,G>eو���F\���[̃��\�C?8Z�����u���
yD�f��y谷/#�#,�X����XY]ae�,--H�M�'�h�?hI�B��" o)�&��e%1�AF@��a����� ?)�'l�%k��:����ɺ�:��g�^q@��5�|��h�i��944̌�8(H�OC���G�<c�s�y�
ŋ����凧�������͡]�<�q8<-�~�Lh�,��z]0���������������h����y�k���_Dr*��<H�_����219�ˌ�T�|�:�Vy��/�O��2��{�z� K&�}�}D�h됍I�%�V������t�	mlR/N��e�\_2�y"��ڋ���k��u�,�f9z{�ࢼ~#�{��;:���b�Ar�.p[1ȷ�z�!hl:Y�S���~�!~����[��^VWW=:>>��#��q˼`��Q=��J�4u6U�} ��d�� ������ese���q�ezB��p2�9���Z��Z{�C�ۀ)q�����9���-^��@�u�{��I9⩉�8Ө��t�.N��T>�ױ���t뼿0!~b�w�`�O:�|y�vIʗG����Yn���$��ã���������Gl���S�K��	S���� �j��@��
GС��~|����
��-��m�֩\;���f29�A�'ǜ[��2���m^����uc�	�8��N<�>���ѽ�a��*'��r������Ç�$��"���:=��ҽ�4>AR����:��0�e�c%o> F�p�B��%(�q�$���Arh��""0l�Fj1�9���Od,蓦BY�)�#:�V��(�x�J�U���T����(nP�������vO8���l⾫��T���1?7�Q��O�E��˧��K5$�j9��N�����*�"[.��;�4�����ĸP�,�`j���C��V���	�˵�COO�x^����,��ot�Y���vy���� �S'�1��2�C�σ���oz�;�������d����۴���ڀ�)c#����L/����u�J9:�)[�������¿.ےGv���z^�(�v>I�̡?bQ�z�Ұ�1����'�b9���+��/�Z�g#��Su����{�鲲4_�f���T������Z��ܔq�)Ö���iR�`�T�����q�S/�By�X��r���.���s'�܍a��f\\X,c|�
S�J�B�2:�	,r�>c��b��}.D�*�"�r�T�`�[h�Ѯ0m3r��XL�\[n��/{��Uܡt-:����
��<:��܅�+|��X\�O@>�]�?�U�t�^��>��_]q�����t�o��v勪}I[�J��CLqk�[�:Fe�Q�[oT�5e�x�����ęi���,*��i�<� �3@����{:��0!\�|;�颫� �K2'0!�W��1Ap�0
� �B����D�`*�?�?@7�uhүn���X��m��������Q�C�a��%4�ΒG/pfvJ� �7���S��2޸֨+�wC�n��@�;B�1��	�|����yS��X�H���Y��1�N@�����´\x�+1��-Q��ʍ�y�苙Ժ+����1�UύR�SY0�e�K/��|&�;��aV�#S�dLMX^���9񹍸RQa��)1���\���N��")E)M�����16�S#wm%�zc����Uy@��䘷2cU��LO`Z{L+���r%7��FY����G�����ru9)0�}�/[F2/vR�,��a[��m �و��Ƿ�|Y��?������_��$���	x|�d�#�����D-������Е1!)��1|4�d��oOfG����A�{��DȤ|͇�`�i����?��.���#Ktl�'C|�wۇ1��zOF��n�|��c�3ruEFIT]!^�t�%Y�M��Z\c}����1��3^<b)ZÛґL)~՜29>\����\��`\���	��;;���y�2rtr��UM�R
p�O�o�t�:��u$ ��N�en_D����M+�Ke}Zՙ���4��);W��D����#�����1��a��h�8zn�ߐ\o:y��;e�z���;H0r;t���:��L����̤��2�K[��jl�Ŝa�j�ܑ�-�%A~3y �NuD�@�Hnc�1�EA���ͱ����庞`9Qfg�h�y�l�Y$��;1��\��&�F^䯱k�:_�!�l�4�~(����x� �܇ӧq�۞����x����?�ң���Ԃ�U�k�qWO�i�*?"�=��Rj�W_͕;�X����9�B
�3���0 ��{)A��B�㿳���8���
g�P���L�+����ٓJ ��_M�غ�G޺�N��zd�md�@�n%��~�H�y�,\b^�L�cOXU>aqv{�b�ϼ#R�g�]�J>��46ʩ�9��OV�F=��(���'�R��{x|�D����3��3�Ȝۅj��L�{���A0�@]O���#|�����*���r6��N�� ��b��ȍ�ʄ��!l�����7�Ԅ�07�)ZeIy�Ha��h���n�TC��?P	�d��G�e��\�&Rv �q+#C���^��ً���g�Gv�ผ]^{�������R��?}S����9�t��h��HQW;��g�P���}}���2j��/�� 0R��$U�f�����ޏ�Ax�������e������?���[*�/.��i�A�)�P^!�N�k�@��������n�D���_>�N�{�T�=��X��;k�+��7;�����@4�+)�����oц-�4e�!eǶFl�����������˿>-������/Oe �+�j�/��X�׍d����\ҡ�q����tT���҉�r/lX��C��y_/������	���BOq+�a
��6Z�����	j����޺HĖy�{�g2je���<��ln�H��E�9E������t�~�/�sF��λ�:X<21�Q�r���{k�}ɣ��O䈏��G���y�%���_�Ɣ�q�$E}D���w�'��zk�(��Ǐw��FIUȎ�'�=����׽�%u&%N�H�`��lo3��@u�Ta0 Yt��/�%r��z�����7�U��6�>o#r��(�M��![LE`����{/�� �ݝg�oLa�F%R�Hw��u���D-2�l+v��rY�Y���u����rKt�C�;`u�{���\��|����P��>���ۂ�Z���*?�탴bkP`{ �O�=~ ��z��5D���It�z�"���}uݺ/#��}�7
��;�kȨ��4����4����>ƥ���5/��Kk�7.�.� NUVobC���1'�QA�zDJ�gZ��ܴ�[N׉�T�1�|�x?j�
���HӰ�[�3@�	�Bh���)T򫊊���'~z�F�Ee��bCoO���ӌs0���-е��Nm,ZqQg�|����%�����H����*�Йј�>�1O
cqkkG�A����rc{*N�bu�l�WcC�P>�($d��Ov�0v��
�LG㏑�8�)��r!�3�����/^��8>UR��j����j؟�'O���~\Fp�P��g�7����|$�{E��K����`�������X��S��6��v�[�8ۊ�F��J
��Dʰ��e��V����b xO\�{~wA�ĥ�dW�E�ҏy�x*��q�wC��秡���3?q����&'�����׿�#�?����u���l��A���.o�Fq]�pè��ڐ�6mʕ���#���9jk�V�i�1j���A�#7Z������/�?~�uy���Â�2��"�ͭ���ӷ���ג9v9��Cސ�6�Fq�m���)0������d�S����%�'��dT�5�.�"��)���sm�ߗ}�oe��ݔ�Ĕ�+:��^�㨗	�^�V�A�Y��}7�p�p��B�]�Hg�/�X_[.3St���8���m����ݑ`KF I�Zy�G`����@a�܆v��p�Ȼ(p�U�z�7L��f�m�f��HK7�x�V2E��x�=�k\�?�=��4e���ђe��<~Gͳ�����(�D>������}�|��[�unM�y�g��G�=��ri�+m`8�
Ov�/�� 
۬n9�A6x�ٻ3��Ň�u��gā0�?*)���1cz?⍷�ؙ�ާ'���a��̡��ܔ?w`6�W�.*����e�Y�4}���MM[0[���9}������rtr!�D
O�X��7V��a:#�WLM`TO�ɆO�/{��H�S:�p(,��Jˮʣ�@�EO4̻���+�޼u��B3��}��o���{K�sn��9�S����I_I�D�||���t*�L�K+}FHl��<=c8\�~���,Ϟ����F���ʔ''���,�/����9n�������-��Э1��1ZC�,�#	�Q��5d��S	���m6�(�0wgO��O� {B����eԿB~�yX��=�;���y�Q
�ǈħB��E��o��ny��Bg�߭0����'���KO��SWh�wU�_�xS���_��Cy��9d�=����FgЉlttG�~"���`���.�6�_z	�����'��H�O�!+�ח�w_=)�|���/ϗ��� ���Iy�j���ë���[o	H��Pþ��W,��B��Zw˰WuE�^����ӣrv|X.ΎU98v���˂\�B���7ү��o��m���F�f��Bc��3�2�L� :�w�_�ʷDC^��-N!�4Uq�U��`��r���V<ݎjF�D��d �o}|�bEƌ��#����T�~�W^D,��=aw+�L��b�3ed~^�?��w�-�)�*�0w,�]�����d�����2/�ͨ�dP��cJ��e�����~���_G�t���
�?�6	�����A"��S8���ݘ�~�?��#?Y&�E���N���jܪwzvvY�G��>�A�ʙ
ª|F����`�K�\���O��d�����D8��0�QP��z��cDy1���b=�9-w����h�<�AF`�v*���� A�|�_Z����r�T^�)��8��ӳ�l8�g(c���9��m�%�Oʝ��5���ݐ~�q1%$VB{�Z��\c��p�3��n��~��9�,h��!z	Z��,�d�2����)<#����<?(����qXyP��
V�(媘�������[4G�1R��*��1J����J�[P�������p9�_�9ҵ��σ����oe�b��N��o����V��Zऔ��Qx�������C#��"o�!꒧Ȁt�+��,Dw����E �`�Xe�2q�9����d��sRWezz���ΗG���G������k�|�q�����{�勭���C�KHYA�a�u��Y���ٕ�+NrV�c41*H;�\y�崮�ҝ��$vG��;����D��<�9�����2JΠ�\�^���#�HZ+����L��~ɩ�|��k#���������eyiA��t����\�v:CGji'h}P�������B����C����@�T>���۵���-�(�ܗ>&���Y��C�bq����N�K1���T*�I�j��i�۟�lG�S�d�׆L��7d�ACu�9���jV{`8�$f����!p������L���w�u�խ}&!����ޯ@�P�V�b#q��;اA�/��2�bK0�2���?Eͳ�-�<�q�kM��\��na��Ť��{��}A	E#cy!��1���c��Ύ������f��e|�DX]Y�����tl��x|B�u�7�y�M>��v5��[�2���5B�FZ�=*E4�Ee;���%�vcˍ6'����]]aa��`��7�~��E	*6E��J���t7��۞�-hq߇��c "G��}�#m7���������!Ceq~B����}��^Y����a>��s������x�	�������~�|jGyi�.��5�����ҙ�A�dd�N�*5�9<�����QE����A�+oÐ��t�o=0	�*�c�n��u��+f
2�;�0&I���q�t�2�ꞣ�9A�8�����e�x�6��:��aTL:���M�uc9��&V���C��1F]�E�u�H�����dyg�g̕����ѵ�~�|��x�F���W�ʍzw��t#��t!��_?@��R����8�A�1�9�1�|�f�;˰>af���d�+'��2��)��w趄/7��֝	��$� �If�rԓ����Wb���#�_u[�Ve��pL�[^]�T4�7�V��]8Y��b�X��V|�����>%P)�!兘{c�����~���g�}{�LMx?���yD�o/��|���t��f�85�9ɬ���.)'+[ui���~�x�Y�5���I���_�e��M�f�X�> I�/1- R7�L�?̥���@~;�yT����Q�P�EaM�.��Q�L��ƙOzT��FnY%�-v,#ll��������g�8L�]���\���&t=w�?�0>���Ao� C��6���iW���^���xA����Ԙ��2z��1�}g32�9�#А��'A���(]�-Y���:��lΕ��9`п�CDJꌽo<�B������dwR��a��^}��	F!n$H*�n�ޯ�����ϕ��?�0r��=�)�������])�s�S�I�uzz���Δ���eEe11�� �q�эK���]�I*�t���7���b�X�0z���=��w22m5n�IÑ67�<���'އ����9�Y��>(_]���E*��	��0�i�#����o�� �{�h���M*�4�L'�v�D�-�5ir�Ձ	��]����ҹ�#}��r%�p����z����~X�<���L�A>謲Rk�z�U޾�)'ǌ��fO�a�Tb�Uz���r�=d������� dԹ��b̮,�{
Ѫtp1��~�ڋ,����u>=�e{��۬C�[P�4z����[�*�	��~��y�>+&�W��c��>��&�%ѹ8/����z���])d��ܨFzK����y�<�7vJw�����w�*��O�.#�����Ҽ�Ɖk�ѐA�е�`�ޓ�����FǫqK\���Ro}<�?��n���)�ͯf�ׁ�no�B�KC��SSq�%a��uM�xN�\P̵B����F]��n%{���=��Q������g���#���sr|&����"W�=
G��V����q���G��B�)6]�����{�Z�l���Onrld����{��3��н.���X��n4��D����D�Ҿ����Ĩ7-/�ɀ��a�gqʒP���f��SoA��y�g��ƕ��<�1�|�)����.��>r��g�*+��%��Ԑ�(���VՋ��-,ʑ��a�vG "!h ��2R�2m\�@��X`��e��Y�/�t�_��'��l]�ݝ#5�{e{����oy���Ԁ��Y� 㖽oq�eS��v����!/�%P%�K}�`��҅�5�2���իl�o�K����]y�O���+��d�ָŠ
���I����鐲vd1~T��Q�Y�-�� !"��E��K��A�:��6\B7 ��r�������Y9r#�@�q� |� �I6l�bD��B�]���
�G���{���V�g/�=�ɰz_&��G��o��yR?\W�z± ���	���/o^o���CE9R�'�-��24�N�0��O��bC����y���:�^��1{���h_/��x�Әڀ8(�� �ecs�ll�c�L�����SU?ppB�+Lg���6-���e��m�-��C�?;�m[WI�����a�6���/>�Gpq�Q�Li����:4�+��k��1�9U/AG���������4t��5-����̣͕>�[�����Ѳ�8��hFo�z�.�Qv��!x/��CݫmW��K����(st��w�p���/���o	7�_*ஸ(Cc}��B�s$�(n��ǀ���@%��N���	@�M��!'�FQb�)L*B?�����L�Y��!����Ȕ��NN�s+���¿���F~+r�����:�`�P1u���}5^�D�?#dC�s�9C���d41W�Q[�ܪ�g�vA�an�c.��i*$��u+�p��܍�^�\!��ɮ����Q���⪆L WNbS~6wg�Ue���{�\�A�|��>{����TXyʩY��"����$V�\��4��~!?V�Ma6�x��RF2Hَ��J��HI�Ŋ^5��Np���ܸۥ���rY^�-ӳ�^W���\(��'���L���8�̻����۔��c�C&ՙ.l����?�n�c�
&�DA���PY�/���Ç���:g�ψ0R�̿e$���u�2-"�se�>����0���/\�_����\��?�C���C��>}v�&�>����끚V���L����~�qjBZl?w`����~�D�`�T�{4GY��[#:Z�ъϼ��H�	������ԭDB�'Y�Jr�	���
��@��jd�΋t��5�ٝ*��2=5\V�g�O�˗_��J}�r���\��w\^�|'ܔ���Ž��0ٹjt&x~�eedE���"5���!_렕Q�Ǐ�%Q|�À=�1�քoE+[L����)����c��!IaLY�`/T�z�._L�2�|0��̲ nff�,�����2Ig�UyDf8���P�t+S�h�0h�Ŕ�h;[��W��+�Y !@޿Lm�o@~B���k��t���[Ö��4��.�v�X0��ea�
�C5$Z���˸=�q{��fW�d�ِ̪����/W�;����/�������Ŵ�O�|_ya��  ���5����)���N��1�>.AX%����!���髨�$���z�A�g�63��T"Ҩj�JM�3����WE)C�#,ą?ȕ�8GU�COcv�lf,Gb~�c6�8�4�EZċ�O��$r��Ͽ�6* �a��8*cB�L���2
/ί˾����C�J�v\�=g'�f��XX&㏄E4z�k%���Y�V*��&�)m#���0���I��j%�#���yo�1u���+��&_��ɸ� �{�ʰ���-,� �'/�Z]��a�`�py���=���d�U��e�j�!�U��6�t�E]�C�~.[x��2���!Ѡt��(wF]'Un�|vx #]���Α�������������rYW^������r~vR.NE��O"���Q^<�Wyc���a�w�*=|�(QG��ߤO込]�*�~ltZ��,�GW�^�?��7���<.'�צ|+�X���o�yR���Iy��VF���i9;���<<��骿��rn8m���Q٫���E^�̐R�*����Q �w��3 �����rS���L��B���O�sD���P�F���i�J�؈3�us���gbk���ӎg���v�j�����Gɇ\��܁�^'�]����G���:�~�9�+�K�����%	D�84��t�t� ��Sv�J����b䨢s/"�/ 2:%��C�1�N���R$�#����2?���6_��a���=ϑ �O6�N�Ow����[��}���	(�*�Ҕ�� ��_y�����H8Ny��	�E�}B��әؖoyY�DF�_��y���I�^�K/���~���~S^���>ì�g��ӒF����	�.4�ɖ ��(Ӡ'h���h,�oj+:?��"���bQ�� ��$0�By�qK��f�K���1n�i�2���s���E��!c�u�����FK�O�AAS�-�'�BN$����g.",?;,�R��~��uL��[�[����Z�T)"D7m�x�����C���'ʳ:.cj1Ǒp�]�vM�r�W�n~��P�<)��W�����ou�_�{hp�x��t�����=.��|
*}�����3���Xu��Z1�Z��=��Y����SU�����6m��!2q7��}$�2D��-�5�.�W	5�0�����ұB��Wm�]<��P������o^럣�PCW��(>�����ݖX-8�=���p��3!g��LC
��M2WI�Gne��I�����ʓ��+9AUBs�Jڇy�utq��(��+�$$C���[&ϳ�=Ag��{���+6(g^�XYZ��rX��-�X=_U
�kә�)4=��KS/.��r��2F��f�~q�+)�a�ch\<�'���}��hh���^�(=�ɲ�>W>\)�������x�C.�����B���l�4$6^�OX�/z+3�0( ���!�܆y��۝���Z��g[���oT�5|�dbyyF��r���G�lyiލ,#a4���@cE����z���Eʼ*n<����~§HV>[i��0k��/h�����C�.�օ�a��2o��%���c����_qפŵ2&wB�����O>ڱ2�A8G�L��%��u6 ��T:"`?ք��Ѡ���v�F�5>�P�3Fk	�q��S�]��6"cj�<y�V�|r�<z��U�,ZE�Ϙ�~x^޼�/ϟ�+Ϟox;-�y�2+��a`�֭��;i��nk��`��g��']Q]�y7Lٺq�E�޿�ZY��Q��x�N���M��ƨ-���W���4Bi�<�le���{u��Z��=�� ��+�u�9�L�c>*G�E���\�`�.G�se�mz�`'��ᗆ����I8�Q�I�K��F�͸���H��)-�ῑ�&:��D� �]+o|�b���)osezz�=�G�����s��vD�$JU�e:#ȕd[�.� ��Т�!����p��n=���!�<�k��/@i�\?tH1��6R�=�&�I��.ު_��R�46�
�ߪ���"�@�`���P��^P��ೋ�-���!�O�^{O�M��d�I~���ad��HȝO��2�ˣ/<�aUʶ�➊{��[�d)����2G��D┞�{L�g�&��ab>��x�S�~2��,�.��G�M<TA���]Z[h\)���m���K¨�=F�X����=c�9�����q/�`K0�8d�F�@� ��J�C������íC�i��.m�����	ă�F~ƥ|�{�	�N8����GŤƧ��}�x�|��^Y\d��`�SN��dƭ��m09͊jlW�Q��_�;F�j��xE�x���D/���@�9��3G����>{#��W�3`��*_|q�|�͓��W�������������\�+�U�(��8r����TL���4Mp����0��ԟ���m�r�_M�ş���t?�*��ks���`P���w��1�fs��D���4�pQ����WV2�p��Q�KW�
<�z�!F�%&��30p\.N%��eee�|����������o���r���cQ/�ޗuT7w�ˋ�����,���H��B7�(�蘲P�Q:���s�KUM��)tV y"�O�R���̎Il��*�e�����I��j�C�9������f^��;8��j�{c|eB_�.F� ,��++�
̟�L3W{�b�o��/Wc�U����A>?�N2�dҖ�;�������I����Ƹ�\[��4#��S��*;)_�����2��n�p�a��z��	U����r#r���%�霝�)S�e���B�>�g*��H|�'�e�&��|���\N= ���E^���ZLw���U#O�K��z��P�'O�n��0��}�o���E9�ƶ4�q���bO��l�)a~P��:��y��cx��D�C���\a�'
�M�߻���.����0nU`���Ό{K�e�g?+]c(ɤ 5�iÖJf^9�i=��[���n��:"o\Q�6n���m��91����0R�d^Y�@,�����'�.�5�t���֏���#��o��Cp{��llr0�A98��'��ӓg�����ѣ���$�7��܄'^���'�-i��w�GD�[�\���x��S+D�9��yyl���Fy�z�l�;���jA�����˗_�+_}��<��>7?��!�L'9S|L!=�C'�:���xQ�����_y$ޮ�>w!H4"�<���z�'w�L}m��|�?�2�P��.�t�:�K����_��`����G�A���
�N�{7�؞�z���;�lm�ͷ_����<y�P�=g�x=9�*[̳}�S��H|%��{�^��)!�g}WA"%����:��t�h�9^��8�pD��Ro�O�q��>W]�)���1Fl���:�����'esk�G�n���",�*��wN/t�E��Ĉ�:q�bne(����~P�ٌ��t-��f�#wjjR��G��-���{�T�������O�5�u��G�v�g�$�E��Na*Z���@��3x���ʌ�hZM���R��l�Z���kL`=���ƭҭ�L
i���+�<��� ��,��,}? :��4��<�Rq�U����ڥA�@[��e;���aܦ�۟�o��oV&��0Q�@%���~L����a���m���y�P����׉�2;+%�0�	��Y%�	F�"�4�פG1� pOE�l���~�>���I��&�0�$�s�TQ�s�m^8��嫷V�qB�g{���ٲ �v�]�~�l�%?()Wp�7����^	m8�gB�'*Yw�UqX��H���A����2ҙ"�TV�ɳmσ�2ng���s�1�0�¨K�DS.��B�H��g���M˭*�����?$�q9I���5�ʋW^Ls�_�'F���Ty��R�����6i��R���[�c@+��d�/;5�0�T(k%r��@Љl�S܌��h�h��U����u��q|*����?���֧wb��B;v���q�Z������U��7�NAQ�d]J/���ty��^���~c�veeI�=��;TX�ta��ǧo��ʛ7�^�ޤ��tlu�3�R62@�ʨi �q�6)�ނ4�n|��ŧ�a���rvz��52r�Z++,Rbjk�x~�a|��)�2�����-�SM?i��+��W��C�k�ם��{���'J�^sbzoRz�O��K�6n1��䄩R��������vY��F�2��Qr�v�T�ӎ�ro%Xe�,��!�\iO��Iz2�]�z�����Y�(�q�c�tLNN��	O3���]&�~�Qn�0�Ҧ�4G�
Q1ۭ����7��Lt�~�}�~��	��<p�S�d#��J:A�ayp{_@A�d܆���[�fD?fHeJ&V�fa~R<w���P( *�]=�
����=>=��t�R=W�%1㕙�RұuR���	p�/�"�b�{�����<O�6�`�-�,V$����;B��(�$*���^6R���,s����]!�U�}Z!X�E���rH��Q���TM� p�۰ŏm�?�����f�Gg�_қ���e{-8FX��'�It}}�.��]�f
�~g�B���ys���tQꁍ����4��n����`T4�ӓ����ś��٫���Vy��V5l0G>/�̔G�W�_��ueuλ*����r��'/��B.�T����/i����[�����X�Lu���-�"S�g����`�Y.��7=�!dF�����<@cJDmX07��G?�X󴌏�HGNJ^�=��������b��QŞ���#{����Ay�bK�Q�n��z ��b��[4�O�Ŕ(V�[�=��R�u0�V��}6���b;��@g���퐌t���Ҍtǒ��Y��V���v_�Ν���3Q��"�q�u>�wzJ0������+��y"C�]{�� �e>�{/����t0p��d؎���:l�vpV8Y�	�g6 �s�H:Fnc��K3�+0h	z��Hi�s����@�����(�ѱ!�רG�1n1ʓ6n�F0��/����L�"O�߇ i���[������a�>�<�u���
Uvb��i	������7�����O�ϵ#���?\3�~z�0���<�Ȩ����F������z�,�D�F8�.M�d�[B��few
��k��]�4w	�H�Hh����8��@(�*u[�t&@.�TdFX�����l����SU��4�X��%�)X�rC 9��y��q�և!�u��?� @�` Ao�ǀp7潮�U׬D�5ع��R��_��r��J_�:���j��癞���+�E�_^�}؉� s\�0~���k�)<�Q���	�yv~#�J����z�9R�_:����߈��d��_��|��s��;T��"�������Ճ������.i�+/��-��"G�QP�Y�D4��J����v1�{P��7��G?vA�}9h���#g)����w���_ˀ��~�3U��4���a!T}� ��<��p�xϽ�4���������m�����J�[؊hs������������+�#��b$�@���n�V�+59��NL��G~��1�2Lh�S�*�s�����.��P�~،V^�S��:����|#�YL�'}>e�6@���iy�����Vަe�sz�)���bS��-�"�Yhٓ[b?4���k>ʇ�[fG�a���qrmepY��N-;�X�K��y�|�g�V̇oQ/B'O#�ν�R�����S����	]��v�+B��ŀ/\8�Na�ON�\n�"���wVN=����k"��5y�G� !�O��-
����{�yӝ�냐�,��_i�@�]��A�.	U�����A��Rc&���~?]?yG���_�|���1��7T��k��ՇҍO+�Ri��Ds�������\ѓ=f���X���CQ��~��PXQ�I���Gl����K$Q��ʽ�;W�h����,�Q^��.�q����3���]!.9���#��G�������i��È'�X�g�	����8?g��z�l��`� �B��v��m��Ո�D���./^��>���0g��[�f9�aՋ������� �o���Kl�ĖH��6=��?U�:.x*�T=��{o����qK~�KqS�;4<��B)��잰Y�?{�F����*��Š���,��/��e�~��C��<b������#����q��C�����}2������?��[�t(�\�u!�H����n��3���*��IB-#�Ӂ��>��&�޾��^1y�.�x��g1��\N���G���×�+�Vv��~�ݗ��/��5v,AO���88�,[G2l�ԡ{���N�����hɑ#�(�ԊI2�5K�:�f�7q��~�+f�ٽ����Z�֚�����#2"���k�l� �`i�eWm��c9�`d����[ړ�S����=�<��t@q3~|$�C�u�x풕�{�ny��Q���+���X8��{�z��B����)���W+y������ճ��B��(�%���̦�<;;�~��_Y���-}ҡ�l��Y\\/oޱkK}k4�1���������Nљ�_�r�&�D��=f������&�y���޽��k���Xs�rҥ\��w�':3��V�Ǥ�u��Hl0�d lO���z�]NԷ�Z�_L��6Ǹl��L���t�z���pcAl'ejz��	_A>��h�j�{�J��:��[߃�
�ۡSA|�ST�뗀�)��12 3���l �	�:�%���<i]�i��M~x��� �0�� ��G��
�X����Zb/XN�z�n)�S�VS*0)�c�.�]^���>E�㙲|͕��<F^��d�e֌W���;��k���1�L�~
CEC)e��O�V��e���ƎgLxe×Ϝ�5��}��t�s�Z�q�]f�b^��*?���,**x;[��-�x`b ��b�u�J��HG��y`�f�J�}��My����� �7Y435������_�s4��ߪA9o��E��S�c�H���I�=�{tt��YtCv8h:^6�Tlcl"�� 2���,{�ｧ�˗��9�g߬h�܎Ea�����on�?��a���������Ց�s��J��Q����?�!�I�������T�-�N��b6�;�����S��g���0)����U�u��axp��'A�k展A�5�A<%���P�4t�����{b��\�:�A|dն�V�ZT#{!����m�Y�����#?��P��;�ˬ'_�{ͦb�٫����_��_zQ~��eְ�6+����D<)(js�#�S�؅�l�mU`��	��*W�퉀���L,�eW�{e{s���n��ߗ�����pl��2�����nYZ��6�l�wx =�H��hp�>d�>��klЃ*�9��5`�ݸi�� W�k���Jv�YVf��_*������}˯\��e	(�(~Lplm�7o������Y[�B���B2�(dceK�0���׺e{p؀ٮ2�y��8�;�#tȐ#����Tv�e��o��r���~����x{��,��	��C����x�؄,(��H��K�� �O��M� �]����?~m���RnѯezW�7�`
�z�k��qiw~��3�Cz*Lʩ�Y1�����o�j���okܯh=ȼ%@��2�t�g0rh�>L��dn[?�e�ȼ�t�~�a�:�I�f7_A�+zC�C�!1��e�K��(y��+3�<��%�Ҳ�[����e}�{��>��.�œ�]��R
J�
��S3�:d+�Bu��$['�
`�*Ok��C0`*�LQ8�J�W�7�[�յͲ!yx�g�*0��ڵ��������`P�2�$|�����G`��5��s�c:�=�t���~ѡ0��	R�yE����]���Ä�K�5X]��{U�:$S~I��Nt�U��0�#m��tPVf�p�R��I�SӑԶ�@0-�Ԅ�M|�Ƙ��a�[�Y�E��=��V>��j��~u�ܿ{�|��)��.]�����X��^�ř���L�Q����ر�cա��u ;�����ֻ�Ve���4���幟���4v�-H�����=~��{@�}}���ߑ�����o�͞d߷������7o���u���R6Ƥ4����{��{����/o˓'<ȭz&T]�tC=d�����Ԣ>4o@x�F�6�O2�r8�^ÅB�=}$K{���9���}�Z�u�j��pѳ���]����Җ�fBNPC!d�����mW}ؗp�E��f0f�՛.&�S��s�S�m��_�'�L�LL�/��-���l����[����iy�J:� �G�����`�q/���A�.t9%v��aTV+�3���/� ߑ�d�B���'̉k(�|�J�@��hlX�����c�bq*��N0�i!���2� �n�<0Ý|J��ٳ�c��+:�����1�z����;-�$m��/�Կ��Z��#d�T����ʃL�P�?�lю�l!���gAЦ�Ua�}�$����t:^�b����p.�\P�6�&�W��\�:J5x:W^�ź�=/K@�]][+�;;j0Gz�ః�r��T��'��1�p��
�|�����3:a�	8C���@9e� �,�#d@߇�d�U�PƄ�Gt�(T�~��&�vee���oxV�@aT�:\(W�^�"?=�k�X�v����/����/�ڨ�V��i�k����Ym������%���9��2k��K6��
%Ő�8������+���Xz��2x�Ǿ��]%���Ճ�:/�2S�^�*eAn�2����bFGR�PD�f�'�)����O�͍����Ry��Ey��?��~���g�2=���܇��@<|x�\������)�%[y��\'�Ǽ��e��ϊM]��2��Q��������B-��:�e�rp�P��ج��B�W5*���̜��^�4�<�����wߪn�+��\�b;�-�������<~�Y~�������˛�+z�U�)��Y[ޜ)x�Y�z�=}e�����s'��|\ˣ1}����dv���[���[��s3�e�Yd)�;�(�W�VŻ���p��Ǹ�Aq�L=�I}�ҫ}����OP4J@���>�b��l���K,�\(�$�)�S���zSƸ#){�]t5^��������R[}NB�E�4�!SIR.�n��P���cK�1��d���6��P������l�l�o�&����	�����a�k��@�&�G�X#}��?��w��7�����������W��3���ɴ�S�i���X>�̗Q�O`�)Ԏ��Gk������&e+��^7f���^︱�I^kj��zB�c>T�(������>D��c?x�֯�Ղ�)��������`�vƏ��``t�I�Q�'~B�d�!M�~W'Fcg{ނ��l�r�z��8?�u��o,x�Z���X4�N�e���1�g�
�I��1���t���׋eyqU�ў;|^;�L���+冔��K���e�VeD�4�����-��)l:���<��f���H`�آ�U��0N)��R��v�������w��f�-m8T��^��X�~�B��Z�F����wUFW��ll�W���T��� ��y�y����( 3N1;�4���5������S2��<����D7HL�:���P��PT�ܟp�Q���t�����7w�w���a����)��V���8,��n�'OV˯�,�'���!nů���9�1�'��LmRi�ko������y�TH��(�' �yS�,�D����=m?�!�֭k���[���k����yepyq��z�V�=Y,o�?�$r �Œ)�G~u'��/x�!'�ǟ�o�4D��h��?���r��pA���Q*G{s��Z�O�T�պƟoPl�V�i�0P �{2`�z�� ��Ի��Q���Pl��'
����a�������*o�bV��)�����g9�'@�� ��n���~{�c��]���t����v�����t��C�Y�H�Z)���d��i��QiRpc���<}[
��:iF����P�����0�԰Q��<���`Ǆ�)[��EQQ��S��E)}���g5�$�A)d0X�Vր���d�H{�J��r�J�7��k}���WŻ���Y\����#����r��g2n߹��9�?Rg�=E��d�*ut�Ȟ�7����%~������D9d&z�,�[.O?/Ϟ��<�S� �IC�{��r��)�W���"�(Uux�U�@g�"�X����kf��~��E�D^p9PdHG��L��$N*����eue��|�T~��Yy�������-�c�����ﾽW~������)7o�*�,��<\c=�y�,v�$(�R$?��x]*Łe+��D��R��;�D�H�Alt����!��j�
U��)���p�g�l�UB�1ް����<���	���5��x�^	������,E��7��o7����It�c����}��z�\���g��=�b�Z6�9��|�%�b�CH�y�cN��˜�F������w�ח�Y;x�N{�ր>��{��fm/KY���)H{��ӥ��ϯʣ�_�W/W��.���(?ꏜ�5/��[��!���R m��.x���B-e�!�X�pd������&�����ͫ^B7Y'aX^�L-��ª?����r��	��aF���h�/;���.�.��(kF�{w��w���;P2OIYG��ti�"L�@@Y��Pj9�Gc����?&cv=�����;��|8��T$C��`F䦯�g,��i���jG6��#��`�u�u�����[>ҭW?P�̦jb�S� =� B�� C�	�k��_���>�2����~��V��Pe������z�n����]F��錎O���q5:�]=�7�`v�!3cg����_�OO�C3
���pQdt��9�I�Գ�[~��Y� h������qO(3(��5�K�+����G�H>^9��*Չ��3da+ Q`I�0LI[�C�U2Jb#�`�Uсd=��EO�FL���^]�*��a�x���P��/��Wqs3<�̕;�������i��ܼ��QF��R��q��A�ɓ>%	O'_rp#.�V^+�8C�Ef~pU�1���A꨼S��H��/�<-�^/zV��E/���	f7.��n���;�n�����ϗ�l�ođ/�b0�6��O��ա؆{�B�t����1l�H�+��Ő||?����A�n�z�
�:�6�X�h|2G�@ͩݾ}��S��㱋��}��n�왔�_X��<�����O���\�H�9�0&:m��MB3s��0��^�˲Ѿc������r|o��ׯJY�s�ζ�(����������5�����|)\ ��lK~�W��[��+��^�|
dpay�;���`l�~�'a����!ϡ5��˟ԟ��	��!�0;	�=�R���]�$�!w�o��W�I�h(���#�嶜^��՛(�#���N#��nL�xܫ���T�&�:iTt� �|���Lr�f�8�~��3�%�����/ڵk��=�r�bZz�� M��é*Π�'D\��v�&�&�����yE��Q���F�	���1Ֆ����J�+utfɩ�d�6|�1��ЊnG�$�`�NT���փCuVt��<815�N���]9�pm�v����_|�:a�p,#g�{����2V�S[���~@u:��H����N�� 7�R�F��ٺZ�{����Ň��c��Y��ݻ7�����9؁-Xȃ�+8L0>H��M�=8v���<��q�]f����a a	�?>Q�����}�f��x�mgg?��U�4ko�q٥�s�p����ԇc�f�.~vUb�Q��"_��cVp8թxX���Y.$-
#
�N�u��plTUB%�Ny����E���'���eqy�l��,~VO��^8W�ݘ.��-%�n��pٛ�#��>�y(!�`1���p��c��@%?2\�A4ҭ߽C�zt�y��zv�]ϰt���gB��ΆL����nW�E� �AZ��'��Ε�����+W�N�����������o6��~yV~������s�Y�#P&F�ٵdL�x���v��!	65�ݗ�����ZÙV��$��ֲ�_�߾�2�{���;Ry��C|l����[��5���~ٗ�_�ˊ�F}�(�L���'��2D��Ln3VT?,�w��-��Q�g���.d�҅rqn�LM��^���QI���	|��!���e���囟����S�q�G�V#@j�˫� �������P��g��������a�v]J-�-{ۺ;VF�/�4*$_��:a@���pM=tZ�g��ý~�3��a��`}WD���6腉G\ن�.�X���X���uC@q�Eb��{��|�'�84�5e@N�I�����j$
�ع�O˝�+�ԝ-�3�]�2M����VK/ ��ñIWiEFG��E�*���$���T���7�h�V�N���d%�����ҁ282��`d���F� _����_Q����l�kS���PBGƓ�H)[0C~E�7)U�=+�3���۹��N.S6�:RuĄcȢ��:�	�p�0K/޽��c���r�����8�̖kW�����R��:����R�ٚLɜW��iB�/nq_��ÄI�����ǣ���hm	�w�]`֝��P|��;]�+k����zy�z9#L(� \�r�ܹ�P�޹�#z���9[^5i0CE]�_H�Q^�Qg{2�)��p!"!��n��Xc�G���{����Jy��my,|�z�,����@�1q�LN�����cy�3S&W����줭�!\��Z60�~#/�}?�́|ۦyڭ-��5�'C�L�C��h��uݪ;�U�B�5=����w\Y�©���U +�-���U7c����r7��G��u����B&G��M~ �����?Q�eMm��۵Zw_��/ߨ]-�{��Ff}�`HNVu4�dv�������iL��m�INGf����f�fn]�Rܽ]�ݹ��̰���ٍ�}R�˻�5��A��r
�0���v��<�Bj�K�{�Si���eS��f�� �1�0^�c��%e�r:R�v��-� ?=����5����^Y[�*ˋ�O�ܐ#�rS�ч�DN�����r�i~
�S�Ǧ�;v.�o+O�5���8�������M�ݥse����?J,���r��[[��4�������_B.ҭ7]�@����wW9Y��]mf���A���� ��V���d�5�.�փ
�8�1\����ƹq���}�DM~u�<O�,o�[�GfqW3фU9T�t 4T^��U+��?ƉJܓ��?*�B���e�xbE1��I���e�81츎k��4ʉ��2I��"#��B���`O5�*RT �Q�+r�-�T2�4f�O��!�:!�(��7%>ƥ���=5�#=���\ʸ����1�� �%�5K(�,\gf�Y=K'd��GDdo��Z�K�\�hN���)n2ψ����qv�*џ�E)�T��-)��g��4������Jr�\���C�9)��Rn�?�a礯c:�Z8ޖ=��ܑdF9��ʛ,�ȕ7�V����Q/�?,��4���/�k��ѓ7��ǯ���:;:�~yy~�ܽu���������2;��Q��2q�#��cF�H���U�cv�5���1(/�6������H��/�v�*/ږ�r~B�����#����_����鹔�Ų��_�ovT�Pvw���H1>�j��5�z����&p�G���滣V�
P�q�YV��a��E��^�F�M��6���`ð�l.�[���7#n��9{oE��b5�m���6t�ޘɞ��'�<D����2�~(͛��'f��
/{)�Pz+���y�"19^��G�����m�#;������]�-??~U~��iy��mY�X/��'Ώq�HS�Җ-l�G��F��}&?3US4��X<�F̼G��Q��(e�y#�޳'��>_Ɩ=�޿}�|��~�u��|h:��]�
���by��uy�v��o�sce|zVy�pJ�>��)�~�~/�%,ᎎ��jXdL���.#�-�6<���H�O8��pK���ƥc/[�#��K�ebl̹��V�~\��w�ܮ�n��C4���+>N������6���%[��,���k��g���� z�}��^�<6ӗI>ZƔ�ٮ�%��)��A�d��P1��@�҇����k�eemS�%�'�=��4!��"��|����2�)�����6o" W_��;ֱ!��ß� ocf����I�7��tB<��]A�2�5�ݾÈ�p���!�d���[�	�{�z}
�ASB��"�H�w�w��l�Ȏ[uO�"�T��p&�9n��9�sP��I����z;&qj���M%�7�A6��/����xX*ւ
Br�w�;0�������?�W�V������e?C�(��>� ��g��s��8��A�)boCR�����7!���A�i/���A�`7�����#O��AjD2���m���aٶ�]�i�*?��q=%_,7����x�A�-��$�X&S�!<�e�f��e�u"�	�5�:#��a���H��9,�ެ�g/˛��~8��?���h�|q�ܽ}�ܻs�\�<[���x��AO��(.E;�Ph�<4(q�J��2�T�ty�z�2�GJ�QGdk��3k�ڷqշseI���+R�ߖ_����x�LҶ���쯁Y��R��uP�rK�&��W�ƅ��F��T>���}�_�:'�O�]ΰĀ̂�������.������\�[����gs�	���
A(���'ig�Z������jV��f��b&m� mA���O��� �H�f��|�Q���(O_���>��=��n����Q)�#zxt��7�Y��R�+�h��?�7�쵯�܋[�sz�g�IU�E;��t�eW׮��7�z��<���u��Rn߮������eI�DL�*"�5�n$s�%!�Q.<��X�6|u@�p��rE����	�=)�GR�'���	���,���1鰔��#)�������L�ۼiS}Ȫ]���p�K�ZeF%7 )Ө}�A��J4����')�,���/�.����W�H�))�L(�Үo��޸�V2N�S����P��J������i
��e������_䕝���/\3еw!��b����/ҫA��	��Y��P��[��[�M�M�n�t���0�S�ͳQu+�N������Sf{�c@U�]ɹ�r��P�m���~������	�t��5��u��T�
�`-ys:�¹��=���4���H��C����������']֌��3Qn���Y��Cf��X���V�����n*�X�'��?(B����؄K�jD�%Q�F%�ywr��a���z(y<)��MH�����8��Y6?�)��j�O"��g���C�a@����o B�a4�:�$���:�����ry�j�,.��Y�Tt�o���a���¬(����rt��p�O��!e��u/�_M>�&�u�Ǯ|��~AFz�@����~Les�lnh�]-?��������������-��ۆ-/���g�3�ۺOo��G�8��
k����C�xի��}d�.]�g���4T�{���-M���jN>�p�_$\IG��}?fAղD1:ƈ!��M�1꽔�,���G;R"82�z��~]����������y��̜�o�����	N�R�!�zo�X
TӪ�;��X�͇�Fu5�ooxHT�H1���E��_�CK6�?<d_���ef�%W3e�����DWl����<.��{>��Y@�H/EP�D��@�]4��:�m�~�^�n%H�޺���p��n��=��-�;r<(S�#���K�ƍ !@޿�2Wl �A`oW���aY\�(+����A��N����ɒ��A���|'�f�2؎�x;R���8����(�a�4?_�f�q�b��qrm��w+�T���R��͛��z3R4��X�(K*_,�������l	�f�'$����SWҞ�#А��0zhf��|����ER!S�D���� :�Pl�{`
�D�TȂ7�f;��pJ�^�hL�'��:4�k+O�^���q�A�[v'w}��q!�����׾[R��nꐙ[���'�\�r���ͨ3�"�j�B����k/��|q�Q�'��T��*l�Lc���{Ȫ�<Ah�_��l�N
T:|�/\����E���2�0TV�O"��mS��1��'&��wk����ލ.����R7�n"�p�URg����}_�d_�w^��������ry~�3�w�\�\���2r����.Uz.?�I<9���"�i�L�S�[���7*��5��ٖ.��|��]��g�����߅?��Iy��yy�f��l�ǎ���k��w9r��C����!p��Cd�?\�ծ;�?:�0`�͒��gN���o6�qS��> L���v]o��1������1��V����*?��E��??+U�|�襷a�c%va=9\�K/'⵼�!�&�s��G��E�pM���[�>^���y�a���;����~8�rU}�u�ezX��I��>�g�H���������Za[)&5�`�C#X��i��A��v��q0Яƫm�3&������q��})��ʅ�io��}z���{�dk�-�����=$/-�{Os��&$��2T��n٤ǎk��B�*��|�5 iU�6�qO��-�ߺM��\Y�t�3�3u;G��1ӎr��,�ۦ?�����C3�C��Azw��
�X�'��<��fl��ڄsXA�n�@��D��%�
�pPb�Q>#�.(�e���ߟ�v�)���wDƥ��3�����g@0���ӊ0� S�~+=U�F�K@��̙*)�3�g���0R��&�x�`{gOJ_��y���
�=��Q��K��&�;�A����#fA�)��%:���uV�H3x�?0T�A�HOJ`�����Rn�<�I��k�8�0ʒ�~~�\�1W��c�D�\�Q\�y��܎�����5Θ�d{�G!k�)�eׯ�F�{�B��˥v�Q~2�O�t`�a�����/^���^�>�;^w69��`v�\�:U��]�׮_,�s�qX��M����o9,���@0p] ��h{*��4&8h�^��Dp���(��x�͍mm��?�������g�?�*������u´qE3O2�*�W���u��_��.����P_�����������I�NŖoγtFa���}D_>{]~��I��o���GO��o\��i��"E�NeG��qe4�Ҵ�68���L��A��0���A�X���rc��i���Pli�W���ޭr��M)�3ej��q���^)�k��7��ӧ�|�3Լ�s�Tz~���>����M��|��=����e`W^�[�ĉ�������+W.�;wn��wn�K�/���i��,�;.�;�C�Ų���1͊:�a��}Pj��E�2@��#��/�;�6��eG9���r��f(�Vn�Yrq�\��P�/�z�E'���e��d�������Z�Dkl�1��I��� �\�;�{��^.����V$�b�G�hÃ�_�r:�N�� "U�-�j4�f�}}��\Cz1;Ĭ@á+|��S�G}j��Ss�=���,pBՆ�i�}|0�fj8�ec3��0{{�S�<�FG��8]�Q���}V�	JO��p��D����l�fB��� ����Pi����Q����!\/� ���R�U)�.N��[��{�ۉ�I�}��E��\�1�X>p�Su3�~�ȝe^o{��w��Q�)p���L0��ZbvXZ�G-�z�{��%&��Ka�0;^nh��s�j�{�z�v�db�KK����m��G�����d�t� ~#d��B?����D3s|��,=�l�o��e� }+|S����چ���S���!^�����j����|6n'hY?	������}m��W�q���q�9 ska��|ru�C\Pl=;2.��\�ZJ}��p�����-)R(�~{e�X}��z�ć��(1��/��Z����\ǿ��m^ͰQlϡ�R�Rtt�6���V�@]�qي-��ݽw]J�t��lRn�aie�<�b�޼O��.�˛~��o�� ^��N^`���a2��|7(y��ƯQ�[�~8T_v�\�|�ܸ�����1)�33z8f	��H�8K+�.�y��Qy�F�g�55�G�]3�!l�|���<�}n�%�f��-��P�''�|håK�r3�e�	3ӌ˼udן��=��=H,O=�jP����,H�l0�/�5�Ǟ���W�5�� a��>BTF��Ll3[R
��g�4�}�s��;�
iG��=	f��U�je��=\���jDA��y�x��U����$kuX[z�O���F�[Y�R�J��h��wNJ-�]��{�L�Ny��Ӣ ��+M���+��37�O������qţo��'fZ9Jrg���8D�E6|�xU>�`_�����;�@�_�2�R�8��\ۑ�	šc��#�W-G�3}��jʓp���"l��ԋ�cCr֫��X��O_���ȳ�W��iV4f����������jл)��4�/���eo{[2Q/$�"�����v��H��I�z�vׯ���),�3�^+-;|1���6�ԗ�<p���vc�fE��G�w�m�DH*[�y�R��*V��so�j��A�Y݂���ewQᢋ�kEaĊ�����ؤ��y��H��#Ni��@CD���%9[XA9�sE�4�]&
�COvD�քuwfkQlYGϚTfmQdQj��o�?��C-'1�J9�o����ߕ��˓����<z�B�{�+Ԟx�TZV�<�J戇l]������O!�/�Y(��K�g����N��[7��{wo�ׯ�����2i�GV��o�a�jy��Z�y#}�t�Fٚ%Ѥ7S!��"l�Ob�5���섫�	U���ߗc��g��|9y�6.G٭B����C����b�v}cݳ��k���| ��#vˠ����m��L���+�T�̮@�&�:��tsxh`U~�%��_�pB����HFR)+ʍ<�|l35��a��{���fB�g��+-[��8Q�m����ȳ��E!��-oK���0�~	�V���=]n��#�3{�G|����V^�^*�^/{����W>��Ňe׮]6�]�V�^
,�@��u_���^7�������k�SA�a6f��;�Y������Z������ٮ,̖7.I���WC�f�v;>�@
W�^��yQ�D߽��d+`i�"@��D�U���ܕv�VCٽx�Xީ���RX�뵦g&�n�c�9J�%&l���+1/!1a��z����v���c���r��+k�'���f��[�5����$��_(�B��E�'��Dˁ��i~2Vr�~�m2q���d ~0�"�ȿS�6������A3x���{���W �تI���s@��.��FYʬ
��	�2O]��:C�?�� eO�L��aY���	Wƚ��&m�\��0PC��-��3~|Y�^���1��J��&����on[��q��k����u��z�gg�'Oߖ_�*/����<��c��,�@9Be
?"��1�3��I[J;3�G���mTJ;k�oJ��{�F�v�R�03�m�ߗ=�3Q���JY\^/�z ~OƛI!eB��g��1�6y�@{,�,g!�ԏ�/�5Z���Ԃ<��+��^����mZ��-�&r|���S���^��<n#�
_4��K�N��$]��`�AO+��	i�u�濂�т��Id��7�������i�� ���
4 ��u�
Ը��ᾚ_��mA���{*f��]j%����)zg�!��,�3$���Kul�${�N��V�'�����:��H&�!�gΤD�ZH:.�^�/���<�	:aq�N6�4"��kG�Gu�9����ٳ���ӗ�͛E)M��{D3S�|u�ܾ}�\��~������'N۱	i�JۧWYY��̝�"��jA@���*����`*�NU�؈;䜘��2?]��%��[d\\b�u�O�4�\�����+�R�/�K�.�q)�t�|H��T�����K������������v��6�O>���!]��v�S�-��=^���r�ܦwOx�R
��ぅ$��vnn���>|p[J�M�ӳ�y%y'dEسO�\oq�U?TA�����ġ�C a�$#rKy�ILς��D�����i���ؔ8�:��#���7� ����z���y
��P��\��1!�V��M��J�i@�9q������p�؛��ty��`0
��tN An�O����%7��E���u��u8�ա�u���Ǻ�`��@��Ժ����7n������ nNF 24i�����l-߾���S�:�Jw��+��:���
ϝ;*�ӣzh�������a�6؃vk縼yǬ�Fy��my�>�-��h�ci���ġ�J9dY���m�����DsϿd�@���7&Sz�����n����X��ɕ���r���rG
��2˾����-/��Wz�g�^����e�*�z���7�M�ZVc�9�_-�(#��#N\����+� h$�]~
����(�l�v^,|�n	�������k�b��}=�0qĲBvH�7��I��1��}��l�@`ֻ�R}NӬ��1#�t�{5�m�i�C,�p��4�/t_V���=�*}���V?~�ruP.�Ǎ���k�.�b|U��tǭ=5�OJ�Z���~IY��$rɴ��{;	&4���ihҭ���%�u��V����ѿ&T0�0n)��_�O��0�n"@��SM{Ww�
��t�,[�0{���[/Zg=': �'_]��Ųp�B�ѓ4�� �ԓ�����I�@�6Py;��<t�Xy�#
�U��'��>g�s��:�7Kq�ko�;���Ĉ����pjF����v@���ʭ!d�p�ԫqu���]f֟ ���Y����w\�@9dkv�`=1�-��!05�Z��r��By��V�w��g�g�5H(�d��x ����;��A����@d!J�gm���b�KJ�	�+qȎĠ#����� t�a؁F���=eqt���0w �����S>�0T�@��
�}fb�o���	��n���E��W�Lm)���s�%����1U�#��|l龊x��x�ޣ�e���w0��M��~�z�N��V�*���ڑg���}�/���̌��z`�{���e��59)�P�𡬮�_X-O�rt7'�m�H��վ<��ȅ"-��oޔ��?�`�"��g�}K��|�.J�ў��|<6pZ׵��}"�}���k�Ǒ���O��{�����V��r���.�����_�!yt2�U��|�j���Y[d|���G~��i��3���ddd�>�Y�D����h�,���$�I��?d��|��rLH���_d�Ѽu��kWݘM~abI�C�˴�����{D���1��+J[k7d�n���{��j�Bԅ�#aV��B7�n�L�P�� U���e����T�Q�9:%���t~� S�x��C������/�[ҵ������n$�=�΂#jߩ�ؑrK�N������űr�������fbrTx��#�_H(�.�~�ʏ��z�~&H`�RPp�}ay��xE�b���[ɺ�5[l�fP��U�x�+�܅�2.Y��dV��X��=�m�|�������g�É�g�%�뿞�q�`\�8����\_�-ϟ�-����Alm�k�����T^��҄xX~s�K/�)����-�ʐNr}��� j+�*���t�< �;�|���6ϫN1;�,�ڴ䖗��(�'�SQ^d�oӷ٤?+�ѿ�]��8f?�EBO 2�A!H۲PQ&���鐃Ud#D}E ��J������i�6��c���ڝ`�}�=;ؽ�{Et����2��$lWi��~(|�{S��o])��Ƨ�G��h,����P��vʣǯ�/��҆@��q�kSS�:F
'���Dqv�H����D> sbu���=���2}+�����g]Q|��r��h/�[�C���X�{��+���_�w��EE�e��r��/48�6ݞ����]��jE�7P=����nj���u(�9S�C;�ЯŲ���S;'����9+�SӼ��7Tz8��>��C,I ���q�H#C�ruz�q�M=i��[�Y,���hG�,$/zOhG�(�Zg�~�D�Q�aq��]P��Z�dv3/2N��bť}��,��* f��V�*g���ĉ�䅳4$)�d>�F��	7$�:d]�ʲ�5Ny�/�rci��
.�.��{foG�@?�>�WuRM安Ҟ�]$�p�
A3��F���߬aZ^�(�_/J	\�{V�N���C,)��y�:�|����(� *����d��v&�L#a���31T�N�ʉ�B���H#Wl�F�z��6� ����y��d[.�[{�왡���@q�<x_S߹s��_�e&���FNZ��d�<7��U�|eYgkCɭ(�T<�S��!����F��Q�g������p<�W��V�7�vVZ�F����YQ�.�w4i;���S�����.�_׮p�Ժ�r��ĉ6�3�ޒKvpE�IOzv?yO�������I-�7�y�P&�F���sVl�޹^n^_�=m�̷Gz��)o^��gOߖW/�� ��5���l��Z�!�?�G&�dB��bf�u�=�2)[E�qs�]��0�R�`��K�<%�#���yyiӇ�0Q��ZT��Q�ʴ�|J��tֶy:�8��Il�����qRU�M������:k�>ų�S���i���,�c/eۥ�������<Nid�n�]�ۢ�@w�7�K|�H��Ր�k�E�s	H��4��S��zL����F�z�]��h�ӖA[H\�Q�gD1*+zPِ
�g�H��.buB�M�M��_aRI�����(�zG6�G�E�C��61�?��Y)x7o,�[�����Tǧ��}o�Gʭh���� y�&�J�Qt*6�,��b�i���FY��0�48��}U�=U8�ww��jA�]n�Z�w�]/��ΗI>�B�2!:1�&M�V����y�����j�Y
,f��*��(>�����G�������]^�X,�����//ʻ�M���'�]�4Un߾�����N�.e�Pp�����#��2�S�� ��:� ��O�QORFZ��rZ�����q����=s��뮮�t�\0U�<���Wy�����`�.��*3eg$�ph�B8.�[M�w�k@+�d�Q�S�ƭ�G����/�.3�DB���l0{�3�Vns�*
.��Q��\�ග�:?cyE�~[iAU},o&Y�95=^���A�����r��M)H�ʔ��?��}�z�<��Keyq������ �����K(�n��5��ޫ����3�«�&t�3�� ���c�|	�����z�9�f�+���E����e/�b�r���s�M�9^�CMe�K;s��Z	Ď>�
�)�J��`׸��)��Z���O2f2v��ו+�˽{L6�,���ȴ���>K�͛�eeeEn�����h�>�8hH�W���df�(w�q��%����e�2�Y�֛@n��q񚨾~m25�M73�f/���@��|���{	�D����И�kI����<�Kd?
���\�����v�ۥF|�q]�6_nݺ\�Hٛ������	4��H���b:�8��ǄK����-�hy/`y�;ݣ�����emu˯�Pp��Ff{��Q	{�^���`���˝�7���Et���6��s9�̀ s���{�CA�j��Îew��L�������T%��׃�zy��My�����\���, ����@r��L�{�J��������d����Z7��	E�G���Y�b�ָW�}�􀤓�:b(�1���Yg�vx�\��?�����;�lu
�C�!jy	��D��������b�l~��� OgZXyoԟ�1����%S>�	[�L�}�� n �`�7m=�_�h��OÖhԯ�ʬ*��ái��}�ƾti�ܽs������ݷ���k�dor�a�[Y��[��}�~��N�A�Eb�6��J��l-�ȥE��oS]����$t�� i�q)��k�R{���rC���� {b���7keqq�Ǫ��X���,_��!�\�����*_�؛~]�O@s
�v.�$<��5^��c'eơls��k33�1���ܪ�[��e�W,)�$:�.腢N?I��\w>R����� �"9�3�&��	��/q>��OH"?����+ԧ�i�����Y)����h�*_��xzd.��z�9ا��8g���<��o+v�p�(�M�!�\ٕ_t8�NKn��ѡ��X�DGpN���������81�]�r:
����=Q_�V3t�<ez_�ډ�ڶ!�W�a֎ �}����1�f�sB��U�|eʶ`#���z��_I�/�g�s:���|q�9 a���[d�GBz�Z�E��ǰ���
ò$���#&k�Ŀ��I&|��x|r��ʏ�3�7���m������'��9���oy�l�Yb±�ׯΖ�����p_�raV�Ǉ�r��Uv�$ہ�[����EŮ�M}��H
_I��Wd2S�k����]2=gX��K�ux���X���!�LF�Ra�����3h��8�����i��f@H���Gw�n~,�J��+M]M�'��W� ��A�� �N���ͷ�ZG�Q&�ݿ���t@����0ԟ/��̶���s�7��,�A&R͘���
��S#����O��|���2?7�k��Lw�˻ŭ�˯/ʯ�^x�@�+����j��)9~��+n�Kޟ'��t�Ҏ\�OJDF!o�&�G���w��ݻu�\��P�ז1���|���F�X��=�٣e|��#8j8vȢtʵr?_�䦗�:f
�"��_�7�����D���FyߨG���^�ׯ_�8#9o,�I��@B�U)���S��o�5���nEZi�a�+Vpuì�m0ܹR�ջ�O�I�ֽ��@�l�J��HA)���
ȑ$� �hL�Ɠ���%�L咉Cu���Z:fs�I��/�t�(z�Q�n^�^�Z�?�@$�HX
R��3�q	*o�� Lu@����\1這a@$��5���c�Ї�e5���uu��N���Yf����y���Yw��!�瞹�e	+�l�!�n^�	��#\�q���.�����'��g���Rd��Њ�/��ǯ���+dkTggFˍ�s�έ�z��c��2.y�خ�NfPI+>*Qd�u/g]�:@}�:Q��FВ�e�ܷq��W����	�{�7�˗�
��W�|�A��S��]�0Wܻ^���ܺ������5X�ܥ��(���?�v��߻e.0���L��\���Q^�o n
oz@&\�!�������X$�֤5}0��zԤ�D�W-�${����]�C#Z�1=NhaWf7͞ ��9�����k��*�ƞr���tu0���i_�q��ܛz˭;�ib��D��V}�g�S݋��^X��=Ч�߹��������q=�Ϋ��*�=�[�ݾQ�.p��ڮ��v~s���b������qvN�_�`R���'77M�ꇆ�-SH祔���JWQ�?�]{�O^�������r���I�ʕ�����ƙXN��������%)�+[^F�=�l�r��?�m����J��>]�W�ɼэ� �H�;�-J(&cQ�%��-~�I��٩r��B�)%�ʂ��$����ɶ����c�%�М��HrI�%-�"�H�� �U��bqAa�\5���!_���#u���Ş�LK�o���a�/M�Y'ɼo����?��0��:�6'P�hr��%횾)8�Ԯ�3 �i�9�Wd0Of��I(���*NF�hF"<&`3�Lσ*OI2SY��1#�JF� �X@>�#x�	��#h$�,�ҩ�CHq�l�HH�N����[�F�`�Z�'&�"`��JcTO��edlZ$G���q�(^��eM,��8'喽`ϕ�_�)���eŎ��B9�$e�=r:A�AG&�lD�'�Ry����'��Vt@��B�
��	�y�2"����_���Ͽ���展��QV�x��X�s}�<dy­�~�_�������c'q�N˧�PO�b���_���-\ԡy�Yfx���m�sT^s鞏�bi	���^v@�c�� ǧt?R�������ɳ��vi�ln^*��Ӓ�'�ʭk5P^/�?�]n�{B9,{�kewsMJ�˖�w8�Ss�\#Z�*'�����O/�O>Ynm��|q�����=5����5�m���#fC��|t{Q�Q���dȄ�(���� k1����n�J7�Y�,�H5�]���;u�AX���������g�nV��m���D��45��B9̫!���χ�^`�5]*�'�]�3����}(�N9��Dy
]���Y�CRP^��X���T7Ω���k� ~Ա��vz̶]Y_s�Ta����O��.�6/C`r�P}�Q�8;Z��Y(���N����7wo�Ks��7�/��R��.픿��y��//����ؑVLcR��+W�K(Rn�:VE�D�t��<�t�{����n�F�Ǩ�;�� �4e<	�I^�K�+R��ɜ*ׯ]��~S
�25��x�lԸ$��뷛eyu����>4�'#���.#�ݪ���9VY��3��7�]c���`/�[<����/{ �9�l��(�($?��y����T�v�Jy���*ǙN�}�>Pv���/o��ׯ7���H�����2����o[9��g~s�4�aٍ��7�HHخi��	ԟiy��d������j	�Ӥ��*�]E7�M�:m$ۭ�[i����e�{L�ȟ0��dA3���	����*��9y)��"�PJ۲�:d�� ���TS��si��P�HBNLK�n�&~�׉�� ߉�������{ņo�n�d�6��?�~�#���k���BSD�M.�����fx��JG+e�����ۨ7�����Z&����D��M��8?�L�8_ݒ�+����ҏV��}���Vû���3n�Fz�1(en t���c_@�zՑ�3d�%��VPp��|���"��x�~x��v����"���N3��0�0����f���dm�@z��9���1�Zn�[�-N�a��t�{��9=J��\?���\Ϟ�+ϟK�}���T'$�v�L�<']�/�^+�^����|²WU��y�
�uŧ;@ M��ȋ���tc&�G;���*���G�@�N7m%�
խAUbP
�@��E� ����tQ�&�a�N��`�8JGfC?���oO@��`u� ��B�}
~	t��k��}�(��u����jQ*�.�T~:%����Z�P��u�z�uU6�ASq���Ed�ſ�U*�(�~}�n5�jevj���)�������r���23�~[1XR���͌��o�1)[�&J��������6���-�@A��~`��f$%���j7��a�i��v0���LVH���{�Ur�?�UW�\��WʕK�~�J�y��]^�^w_�A,/;?R�!�J�� +1�Ee�#��wYs�,�Of�$�7���ޙ'�t���x -�I0A�[�{��X��Z[fm�^�\�&U�2����Fy�bE�zِ�la�r:��d��*<rFZ1����_�w2 �˄�EU����
Sӵ�'嵝�N:���k�}S�B�˶n��H<��+����=�!څ�Q霄�?��{A�~��@�q[��T��x}2�Ȕ^�̫̍�m�>-�R�]\�]�#���k((���ƒ�>�� n��"FB�k�jܐE�6x: +U��g�v��WV6����rR�$J�u�����F��h��`��u����,hŮ��w�KtP���cⓓw|Q*�M��Գ�/��ze��W�zZ^.{z�7=��h]�8�����2!���i����{��A��$�4?� ¼p=���lU���$#3�<� �$_H����g>vsqi�l�|PYQ�(���n�X(�i����+?���_b��~���b�g\���8��ё�%H�:{�H2�B���4��c �b,MP���d���%�J�A��>	T���	T�8W-T�0	��q�%�W��d�Ie�u!��D'L_���p��dU�,�)��LH�	̦6�7v�0>���¸NB��\(��&XR\]~ T#�ӣxxB�ٝ歌�C�S�%�����!t��o�6�K�SRh��������?�bk,�CE��?(>^�?���_������©�|$˰3�v;1=�>�m��Iڼ�F{'��y�r����-t�H~�&D��)Vhy��8�ZH�e�A���=��VH���T�:_._�/s�3��	�C98�P�7y���r
#[2#�rfjysĄFpg���6|�R�b8��U�(��6@��(�F��]� 均��價Q�i{EJ�e����c�mgg�;�<~���my@�{ң,�'�z��D�jx!g��pqߘ�Qk~�y��\(�2�,�	ՁH����3�lU��o0|9�.0�|<|��
�%
�^Y(�J6 �w�-Q�"'�[J2��~6�	ۘN���߃u��1���Çe���7�����W=PQ�.׮^�^��⪏-Ǉ~-����4d�+'�[�V<��9�^Q@Z���,��VU8c� ��ǌ5�-/��i`c�*���[|ԡ�f|,fo���6v��X����$'Y�UG�ʭ�H��|����Ȯ��)^�3m�;�dc5KL8�rC���X��3�(���l������1�6W>�Q�������m�y�g�]����,�LFC�V1�L�3����م��G�>	�H�;����zP�J�-K;)Z�_ϔ���}���P3신���>%����A�l���Ȅ}��������#���W~M�I�H��+]��oK�ۖx�e`W�\������o��C;����յ����j�����_�K)B�������;2v^�-��JB��,JqW1kf�����ؑv��ꂥAF�QZV��[�� 9�ƫ��b����t�q���V�/���m ������eqy'�B�xSVV6
�����954u�c6:���}�����oʐ�����Jh�o��xX����7*,A������8.�|9b<�x�`R���w�嫷^�8�{�I�1�\7N���Y�l�D��BV�UH��}�i�����A�������s�'#�
к~C����Zgkwɵ_1��1�Ua�p�6�o�N >]��Vx�I]��JAO��$e�鏒8���7�f{���#7@�j�xq�\�>���5aT�ۛ�K�c?��T#�:���K�~��Ƽ���rE��x���A��h#>��ϛ7K��vw��K�紟���`&˭[���^`�����>�m(�'�s���	�	Qt���P�1dd�i_��Y������DC�g����Xv������ߞ�GRr��8���Yf"���T�{w��Q����}�������qo[��ZwG�=J��<J�b��(#Q@�4ES�N���?
"���p�a��S\c�L���A�����zyVSf[��u�Y�2N����c*��k���ةr�b�q��!
m�x3���e>��� :�R������mK�9_⡚���Se\핾�չ��W6ʳ�����oʯ��P�Nm^��d��$�Œ�m��NJ���F��Jm{ܵ�~��,��!�H`ލ2�6�D�W������k�C���.͗۷o����ܻ{��H�e�3��[���C){�z8W^K�����	��y=>��Y�U�v�K.�@�=ٿ�{̾ʪ�l�y*a� ��0���-����Jߺy�ܒi~�ǣS�s����2�J+eiyUc.��1Y��,-aiX�u�f[Oa�4φ��r�3_�Ol���7rqU�	��e8��/'��2D�D���
4�bjn�!`&�u��@�%4�����y�fm%EQ���ڗ��b������I����2?���͕�i���P��]����������b�IJ�?䨯ǐ-x�b�a)��F��=��el����M�|�M�	)�.L��ץ��\�Ѽ33,i�ko�iG��,���s,;)�]8D��t�F�[ob���xe���d�V9.�_=/����<�X�6����g8����[��Ç�ʷ��� s�.��c�=<ള�i���'�d�|�s^?��i�	7�n���_
�a���~t��B�o�(�,wӑ��a`�y昡Ȃ�V��!8�	N�Q̇�l�W���\R{�w�z���;����Rp�Hٝ�l&_��/^Y�-/�����<�{�潮��1�ߓ���C�YJ����{����2Jm|��}WX����-A���G!� �!fkc�-�1Kb����Ν[囇��w/K�&&�L�P|nlI�}�^�?_,o�,��!��e9W���y��"O�b�!YgZ�똢�A��6��P�ﶅ�!2�`�VK�T�k̈e��^Y�\fU�������w��P��m��U�0c+d3�,������I�ק��f�c`���Ч�v���NFtM�0��q�����o̠ł�l\�>gpd��<qJq�p��R�N��'d&�[Ǭ�M:T����R|d�)����ȡUs�(YHr!������$Dv^��� �����4={��XF:��-!x��f{o��^cu0)�Ǔ.n��ٞ�S:$�xF�X�ǈ;�i5��)�m���C5Ɲݣ�����D;��z5�Q�qY@���3����7�j�� չ�G:"��?�H�����-�s��e����|�]��;3;�.�Hf�.��)��	I����S�e��:��Rg����<	���H7oeH�<�/�W���$��>1� �Ɂ�/�I���������#�؍:�l��fO�Ё#���#��*Ʊ�� ܗ�bK]H9�>��=�T��{����@��GZ�k ��i�{�D�3⃢a����N�<|�G�oo{=ND���~����~!+��d��&5̽�ã?-0�ӯk7D��uK�~!��U�KH�@��A��}���d��<6PF9�I_W��~�b;%��f�o�����l�}Pn\��W،�(w[�A]-??zS��ק���7emU
���1��t��c%����J�O���.f�Լq����8ն��O�m�D����ڪ�`&?^�K^&�����2==��k�O����w�z����i�TC������z���?��Yy��m��9�4U&��,'���91c*>���t����|w��l:h7A|���|�ȏ��eg>�;:ږ�~��lܽ{�|��=o/9��bs&�غ��ӷ��G/����b���DU�oE6�im�]�� �r	�țǓ��y�+�y��z�>�~�s�j�)�DǕ��>?L1.�xy�x#z*�x"t�	�
A���C�d5�J���?�,1y�4[��h�T9�Eۤ�F����,(����M��~Y;�%6z�a���s����E)�?�/��+�hb�UְSiaF�������-������+/�Vd��M���\C�S!�����f�34�X#��S�r���a3i�������G;)��r�..8:�]V�����?R�q�������)����Ӳ����3;;��$|gG
�?^�3A�ѡoSn5�+�V(��0�t*q)n�ϴxv97�x���Hf��H���.f2�K��2;;-�	�[ �ʠ��k���ݑ����/2�����Ihd� �kk���31�[ ?��"|A�k�Ր�
�������0799�(��M(�����C+�l��8�)�:��)Xۂw�7 ;�ر��`�a��|5�� ���X�ގ?��.�tAސO��u�z��(`[C bͣW�nL��5j��~���u�.�a�f�?y�_O��i<#�=���w���6��ӟ�@5+�J��8��6ֳ���o�8X��������w}��܌�&��q�Ρ����_	_�Ǐ_�d½}�m��Vl=&� 핱$� +@Կ'��H����̪ye�!����9r���@ ��u�r�������o�eR}악����m+��ܿ#�`�G{w��,.�GOޕ��#�E�����31Ų�ɐ�
4t�\(f��|�5`�b̰����M�*s�&8Lw���+c��
���!����ʝ2;3Vn߾���[*�;���Kގ��7Ե��u>$[.O��-Ϟ���˞��%|�j لi��~'��
=7	'�%̎���i�B�I*����"�NX��|�q֑Ļ��ֶ��l=I�#�`	�TdEȪ�~��ǚ�x����[�i�*-�c�JLѳrK�M܂�:��.��F��g)��/͖�Ks��e)�7��Z��=�w�I�M�`̐�\$�D��r�W �UA�2et����xT�:�%#�e����!Qrɬ�C	4��R����V*�KZN�5�.��ٵp]Q Eu�.:� $���B�BOg5{�x������`g���d��R�}x?"%���Uw�����h��"iq��W4���O<w�xW���������n���_��T�2�+dG�]�Vi�����o�B(r�D9	l|L�߸��1ٙ	��)Np��kp
Zn�|�9�� �������Վ�m���H޳�6B�V��P�g���4[ꈲ򏵶$�L5KT�UU'� +�v������i'���{(v�Fv�$�3Ӕ=ʿ�~�P]<��6`��VK�mm*��w���x&t�s��M�t���,-:�]~]$��Жӟ�
�1d�f�ƽ���A0�E;L{��t��[��,�����䈽(�+�ȃz3��_�)�q{�F@��6���}��1��-�(��b���c���������U�d� �3s���f���7����嗟_�ŷ�{ ��Xp[WB~=��*��A>�e���a�
��q��2�qO =%u��
"e����R@V��#����O�J�07Y�߻U���A�������P�DG�KY]�b�x����g�?��Qy�jQ�����1)�3�����	�?Ŭ&����]����i��-oH���7F�G��52�ҋ�9�R�}/�z��v���m{��AR�,�XY�)����my�z�l�*�X�v^�"��H�F�g�\��J�x�Z��D.�Эc7�NO�؛,K~lV;��Qli�M�����UՉ�Q��!�o��!S�W�"�)Ёc|Cw8G����*��[�OO����[萌� 퍀��t®�c=�4M�G�e�P�R��'�!�#��Č&'#�-Lu��A�ӏ��<D(��g+��o�EPC����H&�w) ��p�ҥV�`���'�Qu̝/���Hz����	{��"�&p�떔�}W����2?7Q�.�z�&����B��FCL	H7+D�o��7]�i5`׭��H��T��T�3����2��@��)���۝���ni�<�3�ݩr4/�GC^�8�A�:)։��^�ӓl".Y��oV����H*&T�`*�]�n�>��x�25^��><8�Y2p��m�ùGO^�_��,/�.�����1�*fry5z��u�7�*���K~*e�� <�f�P!��c����d���)I��ђ_�'uLH=��1����d��b�t���?*����w��y0�ܓ�����.�k����{���AG�m�'N�g9RfX�S���o�b�e��m�������r�����7w�Ζ=_y[ƃ:��o�7o6���r���;����'�G����|$ʵg�t�^�<y�� �W]�*���������)�=����N�`�Cp��#�5=K/���lGA�ʌ�eK�ۜ�u�B����rE+��R�������W{�����ߪ*x�C]��<���3���F�R�	�f�.؍���}@Y�9۩�!$�߳��L���`ox�/Yy�a�V���=>�>���巠���E�S�(��V���w�(3�m�>쇮L�X!�6���/�}����H=��z�GO:d"n�*L 9�?Ӭ�6����^6����I8���'�[��l�����kn�TF	�ͮ��hU��FeBMDUv���ܤC5��4h����� 5��
���'�����D����_�ґ���@��2&x����;
z�jȼ� �+ ������8��ی(8��1�5Z4��K������;"?e��S�+��q���3�y��4�'�kC(��H�Ld�"���Nb^�
��;�p��"*@���amF�t��fv��2���+SS�[�+��͍��#TJٔ�˶[�O�'y����M���n�� ^f]W���F�Qna� ��	���6�lc}ztx��}��������V�+ق 3.|��?��/;�{*g�"ARN��"�r�໋�$3�9��8z=�
C�w��}�Y�}W�
�KS��$%ud��P�6������iV�	@��\,��[��7b�Y�q�a�}p"��=��<?;���
=r���R���mm�|���:A��]J�b�{�h��/]�bˉU?������01>�(@����V���E�A}��++��;z =�2��|�ܪ��+�|��$�M���g�K��x;�����*iƲ�Ã����T�d2�Ŗf���� �ve���2n�[*ʳ�+�������t�i|r�K����.�wb %l��_I� \�U6�G�pї�<�ya���f���V�P���[�mi�8�x9�5�?��n��_�xJ,v�Y_���]+��Ų���#�H��?���'ԧD�i�'<S��S�F�>�>H�!�K�Z>�:{�ҽ��ʌ�a4�z��ت�K�ọ�����GІ��1����
��]��6e����Awk��a6��0��:h&O�ת?�&.I���X����6s;5�	��.����5L�+@d�eJ�����̬��d�s�po��+4�ii�~���D*��H���+ U�[^�(�oW��2�����}vv�{������i)Kt��l���o�M�6�V��sʑ��qSgEG���ES诂�O�j��k�"�LZ��*~%���U^�X,�^��^�k������'�k��;7�����9/���+�\��HER��r���aZ�{��������k��,(�L������t��<zY=~]^�]+�*k�Y�ȳ��A�>�K�K��˴!��E�cm�"^9?�����G�T��.~<��M�.������ n�a�~!�	�����"K�P����=>��+.^P��x��[�w�CV��z�v���hI
{V�-o^���mg&vb�W��7���������eҦ_@9l���;�E��`��Ev��W:�L{����e�u~n:N"�� @}
�¶�9� !vX��!B���oYK����$��S:�3�2niPr�����`����k�*t�]�P!���z$�Ɗ�⭾.KѹvM�`�/̔qN�屷{�c�yPY��[B��11&���[�P���e��N�0]��K�π,c�@��L��(����Sl�_b&���{%R����7 p)	�炕�߈L_Q>]�f����7��pkMqR*qe�
���M���n8�3_�����+���L�Ɇ�,Ix�j��.�l���r�FH<?��J
�ի��K�Vn������{f�`uT��M�,�?G��00P������ M����Q��	��)�G���α��z�z��y����3��E�ē�5=�ݹqMx�\�x������ڼ���+p=��mg��^}+ ����P�D����
��a�O�G|�'O���L�H�GU����ϖ7��_��ܯ:_�ZUy(n)���T����r�n9;7�2���wS��G�{�
֌]֍	i���a��;��-������`��g�/0����u��)0�~�&�L����S1��=.ٕ�n��G��N�p0��FW��4�s3�������k���o���=�b�W?^-?��e��o���We{C
�Na��f���L��XS�M��HG��ʫ|�OBk���_V�T@�*� p�70�)=��g�.�?��曞�E���d��#ɻ}(%Eo�li��3�㓓q�o�+����_����޹B�,�v���׊��Y�4qk�H%��w\����L�%y�@�簊��Q?l��E���_�x]�X~�Ɏtѡ�"_��A9'cN^e�s5�:�G��(�i���]?�D�ܟt��} ��̿Pb��1�͘��t�뉓0�m�s:���ځ�|�	=�lE.P�a'�G��$ol<��(���O:u2�&��i���l�6Oӫ�h��-����C=�J��+�.��ߌO��սg=X�<���y�S�Ά6_"ON���E��Э3���?�WSo�D�c���\��:����ZZZ+�;{�T-��x�\�B��Mo�=�A)����So`�L�6
}/-D�f����q �q']�J�fp�@�OFD,�^��Q��9���mlA�_^��2�Ww���I��Nvjz����J�W�2%����;�|��	��f׎�){��\�-���6D�|s�N]���K��1յ����/wv�]�C�_iZ!���cR�fggʌ���x��gL��}�jM��by��My�j٧)� ���0DJ:�;y�m��A&.�/�
y�O_�3v�AӦ�a����n�({���}�0?Wn����N�PK�e���K���9�$ʫ��ʛ�˱���Xn��4�~���O|[(9y,9r�*�dO�������[��b��PI�H��NQ�2I����7�7-o��������x/y�յͲ�w��� 8��!W$ U�~h���y
��B�g��^���"k���)���{%P�
P��v���O�������w�q����=|ĸ汭������`q{����3Ûu1}�S B��v�]F�tm��ٸv %"ls��!U�w��Ŕ{�g��x�d���~�l�5ms'�}"�x|������Y��..�����r(7��鉢'�P�fg�D�_�2?X9��0���F��DC�F!�8߸P�O�Y��PZͮ"BX �4��\0c=a右��-�5�lq���E�>�<5qN�Ty��.les�ד���磫��+���e-�gJ�^y�Ov����#�2�|ͺ[��s��ט�4h��/�����U����O/��ei�l��� ���Oh&oXo,!+$FMR��+gF���f��B'>�����P�س�[<�R�t�K�d���/Ȩ=�;a�k�ƞuLa#_k����B�4�� H&�"QFk
�����Pqr=~C�SP����Q��� �������5�|�Q�av��62�JS�zν�R6�?�wK{~�|���E����U�K\Jk2�Q����O�b��MX�=e]
Jue�����o\��9[� ?���y��x�r�>�׮sH����7��[7��M9ovtx��^�^)������i˞�(|��A_�o�o(�^�)t^��gA��y�}�\�<n���ͼh�rW�����2��;5�%	L~��r��8;')[�ml�����WKV�9(�����*�
K"Z˓7q����P_���f���v������]�#���D��|����
���B�j2A6�h�H�_oA��u��.6�`/��N�Xy�]K�s�R 9� �p*�EҒ���d�E��r���`������
I��P��Ph�🝀�Ɖ���@��Ma�q��Q9�J�~ qj9z�%�"��#/+��f@�A��&�xH}��NY^Y�r�f�F\|���X���"��27��+괏�ݍ{���,_5�!Wwt��1?�^y�:����*�����`��>�ҭ}�KH����C��'��F�$]O.���z��ض�HO��|�{�ܽu�ܾy��W��YF�勳Z?]�̟�g]c���'2m�p��(�z�?�qK����R�1H�-e\�H��>���������������u)�kR����%��e��u�Ĳs���i�c�K��`P�.�F��aH�t�z;��@�G��D~y��j���q����ŏ�����d�@s�� T\ч���[�qү���V�	W�H3E9k⦕n�q�Kds\��a8�p"���i�Dm/���Z����.��ؖ�����[//^,�8�'��ʣ��¥���by���Z����e�F���c�ߋ1�� 8O�~��sLh.�w���Ć��s]�������{�} ��ׯ^.��Vj� ���o�?~[��x[�����2ㆿ���i�rw�[�M��C�?#�CE���O�m9E��BI8���$�+���R�C�AaNhAc��W˭�׼$��M��b�߮�������e~�0�"�ڤi�jO9����.(l�S��~ؙ}ӝ�ՓWNR�af�����eԢ��+��#�Ҁ?��A���n���ٍ��v�P�L�KL��!G����Ŭ|FA:Z/�$N`�D�5�@!S���ȭ?�����O�'Y�V��?�|=���AP�IA7*�꓎B*�C�]i%&�jt2�՘4��#�
3Qy���'x�GD<�[�c�,f��$:�V`�Zp
O<%�.p'�b1��@���%��){B{iV3y11䂬.f\T
����p��3�>��5��!�C*����5Zf9��6����gw�p�WKt2��Yx��Q��/�ՠ��/�:�w�����YQd�g��/+t�I�.VZ�ͧ�Q��0�q?HY��S�ޞgJ3�Y�{x�:���k���+�kOڪ(�Jz�H�Ju��X��B8�$��>�;6h"V��X�RhAy�Ot���a���c�m�x��|Y��/˫7~-��Պ�/p�/g�Kɥs����<~�n��W��\6�ݱw�����]�6�b�x7���>��c�1]�h�Y6iv��k"���h0�p��L�����Z#f~Te����K/f�~�/�̂�#�h��}�I��*�DC��Px�V��1Z��S�=�{��{��`^�8!��'�*��a����e��E��g�,/�m�_��r!�=][�*�����:�
-m��H.��y�%{��>�N�瀖�4�֔t�V,�����Oʋ���X�ό�yv/wo_/����~��ܿ}�kmٻ�谔��Rl���O�_~�xpɻ��	��t��A�v�B=u��O.�£�z�u��+*�ǚ����IqaLwG�_,Ѣ]�ofK����u���w�/n�o��2���_~��7���;��勞���d���ս��ٺ��o�<�2�!=�8�t9�K��L�ݖ�\i�r^k_\����w�:HF+��L��N� ���B�!�\�P	�^��Go��)�ezЊ��.۠��G�_f�Ǉ�+���&~���o��Q�Qw1�%��=�G��%�ٝK����a,�09�6���%X�e���;��JT4��L3ZPlC��F�e��"����V�pV����B�A!(�&ǠA>U�b��KN�Ql�l+̊KEB�?�&<Q`��E�QE�6���{ӱg�-
q3R��ʔ	��Q��<(��ʭ*���h���*׮.��3~�4��f�G�����^��R��S�Yg�j> ��0V��ڛ
C�NG�.!.~�8��[�0�#2�E�%����k�_��%[f�Aq&��c�T�l�Ct:]֩nK�G��q����-語:o�3�?�,6�W�4�����x;2�^K??ʝ:�<�l��ˇ'(���׻�W�R���V�V6�L���z�o� �a[��!еW���/�y���;w�?��;MA�O�1�54��	u�F��R�@:�#>�r1D�~>��~��CT ~V7`hڂ�Fꁸo�����
$Ր?��5���U�~�H{m~��ҿ�} !<��v6sl�$��1D*���8�=d��nï�Wu�%?���T6� _�.����[:�͸и��W�2��F�M
7��@�-�H�Lo�4�J���Gˍ��7����myp��=v���������[?Y*��'^����S�X���MZm��-o	-� �b�P��f+�PVnU>�������]븕@������Rڏ��k�����|��=87;3-����o}=�xW=~S^�|W�w� `Ŗ5��u��T9zdk �>l���tK��:����%.���g3�0��Б���5Ϡ׺���]��z�n�!{"4�ˠ�)<�(	ɛ�x����{Gtz���D��B��Q�>�`wd��u�3!�K8h?�V0�ꭈ����=���D�LM���-�����}nQ,����t̤��|(*�I�E�&é��-�
��C/��E#��8�Br����=P)���ϼ��t*6ʭ�T�J�i`Ǵ�\����OV�У ��G@��8�	[aU:BwTJ_!��,$����a=�D�r%����؀[��}�[Mq|+��(G�9���PE7֤QdT�g�G�	�>Tc�8��G&]�X����qe8>wQ��#�彗V�6\&�'��r6:�ڡ��ǚT:�=)�(�k��egg�DT7G��,�F�*Ny��@����ܛ���|u���=@8�n�ߊ�����I�K�=8*�k�eui���5��,I�]]/[�>���Ɂ��Z���Q���~���<(�i��?;0�,ۉ2�r�z��,�T/SP���1���Ր�pPu�B4�>������!i�zD�Ѥ9�x�
��g�'ɐ}8fb��m!�φ�������b�Ŗ��E96}������a�@�@գ:;k_mخ�7ϲ�Q�r���>�1�@?��j~�|��]+y�=�ĵ��q���G�I��l�������/�ۥ���:�£�n��?��|4�7��i���3�����_�ȋ�M�^]<x<^Z���8f��#v��ȑ���r���~�}m�����~c�x�~�K�����eM�*�-c�S~{ieʼx4
�z xm��/���A�S��-Ԩ�9k�kl]/@���� y�1�zP#����]�%z��uth�L�(3�E���-����r���e��q�r4����Ё�n\����C|s	�a����c�u�7�	ewy`�!����`U��B���r�nUn%�DAto�|�e&r;	N�i���Z4�M�� 趍Æ��Q��P|�.��i8��\;E��X�*3	�Rx���O>6#�ɜ�0��8C�����R��
p��OⵂSu��,£�} ��s���W�@خ	�+�(�c⋏��U���x�<}ƖYK���T�����hY�2Sn߹\>�Y�޻&٧�'<�5y�̅#nuF7���d�.��a���ح�ݲ��U�=�n�h��}�#��_:$wr mH���G���Ao��!���@C�k�A�W���z�+4��oో'�̨���j�i�K��v���vYY^�%�n�;��'2���䋻����d|d�H���q��ᯒ0�q=n(�#�]��ч�X>& 8�eOJ�q�pa�ܼ��Pc��{��Η��;o�Xÿ��]��O}��]Z$���Cbf��T��U���C�}X ����k���l��Z(��;:o��{{Vl9�����>�����E���*�Nv��/�G�^�Rl9����1��ױ���r7��į�n��A2 ��(g���6�C��=��l?v _�)����f��}�`8��8513~ԏ��q��L���3�,g�f*u&��!����%Q+@,fn�ʝ'=��d
-=���[�I�@��	e9�j&Uњʖ�+X0e�UEӒש3��@�[M��s(�P�>gn#���̄��lFg�q��3Nk�04���P<� ��g-Ձ�ŋ��"���''9ME4�o쏫u�����57��������6O�~R�S0��Y�m^�!�W�z�}D�pd�xe�+D��,c�-v�#zJ�)�J��e�c*��� �Hr���I��� �}���%A:^��Q
���I�w��6^@ܛ^�a4^*Cv��:NH"3��*�q�Y/t)7J�;�)�&�6�Ą~�D������mٿ.��?B��u����N`9΢���TP+hoz��{�	���|t��O)Bt�(��=-�Q�"����!��O��W�!!�����g���<K�,/|�oP�L?�}}�ʫh�gL06�wu�Sf�G��[�o�?��;)�7������1���ͷ��ѓ����x$�UYY�.�,��������g�~Ct���!��	U��~������:m�cx�[e��z	���w-�����p�ܽs�|�����ߔ�Wʄ�ʣ�e}�<�R������=/�^-y��X��E%j޻E����b�#f��ʠ(�
}A\Χ #t��F�c惑|P~�g��a ���q-���^�P�73���˹�ߴ�7�r2-��C������-ew<��cj�'>3������H��w�M܄�6�X���o�Ǽ��kW�̭��$��+s$�2�A����Z�(�Ď�ѡ�K�pȰ/��_��5M���/=�g�����^��C�v�4~���\�-wn_.���PwUO�Ӟ����p_�!k��$��]���%u���?j�`A����u���b_d~��uy�����5b��#���X�v}�ܽ{��p�ܺs��_�����e��|��z�I=�,qS�C�9����O�~�x0���3��R�G'���r��1�sDo�;���u�����d��z�����1�Jy���~f
�xJ8��V�?�G��-,[�e�a�*��V��a� 5�(�_�-yOؾ�@���{��*���g<W��M}��/����C��G{e������޿wçW.\�+�S��S�Yw���jy��]y�r�,����F��D_?@��i�� �Qj?����McQ��<�i%jT8�d��L��������k�ϗ���q�]����×u�/^�-o޼+����P2k�a�/��9^q������:b.\�+Vw0�Y� }}iPān�vf��uoo�A�D��>nm��ek�m��~E��2r������y>�/Q��Xu��@hتp�8�����Yҏ����5ww$��@Qf�T���yElEC��-,it �Nt��P���"���@����t���E(��M�u��@�6����q����<t"��3��x���ɉ�����>S&ƥ��	)y��Ӿ�ϕ��=�^���-���8����g��=�Y� ��-�8+X�c
��;��H����~��5�o��� �,E� ��,'����3��A��1��x�z��C;��ߓ�NC�"���'�M��f*K-� <��@�Ԁ�|�软��i���e��3g�<��^7�e&T8��%���&�C�9>f���`�|_Q˺8�<����,�<�g��4;�> ����[���N*�]]w���M0�.�3��?���5}(��^�>�K��K�|�d�v�02�y��R�=��*�'��T�D�$m?� �̗�3�u��W�T�n\�޺{��7��A����������yۯ��I�.3��˗��/}^���3o����X�CZ���S@����8��"�@�څ�O?̷�N<�-�n�bKY��vW���v\�_�T��?��[�]�|�LL��b)��ɓw��_x���5+��ڎON��٭&�Ff����z��@����Ch) t���?eC���r���C�����meL�Θ�@�=1sK��5煐[�;�g�(�@��3�W:`lp�6g޸�_�a?��"�\sK�d�G�p�~�#3�i]s���<�\���n �@�	a�AA(���6��wL���1�WLg<��7�E�
@VZ�S}��?L���p����S>a��Ǌ�����t��������E�RY\^/|D�Q)�s��zb�X�޹Rnݼ\.s,��=�{�9����g��w,�`����
U���|@t�8�mB���f����ˣ����W��⪗`�O�˥KӞ��c�;w�{�I)��Xz��E�>+���K-1���;2� T.2�p";�!����g�c�sq"?��(��Lq�\�=���\$�4?����!p��b����Nt���٠p6�?�9��0*^��l�~pL��C4��`2�K��mN�,�ia6���K�*TA�Ђ�Դ�^����M��O�~��wȋ|�t�8�0�[���q�|�����m�R�(�����LN��kW/�ϻ{�F�qm��L��Tj�����������Zy�mΖ���~������I
�'�󾃩���Y�@��gmaF#O�������y)���<���Eo�y��Xk+R����=�x�!H�މ��z���u�k(y��gYGg0���t���<8��:��g�n�J/�mCa��a��H[Va�Ը5y�
�Z��;��fz����إG�� R~��I��H{�ޘt#�~���O0��dV�'�VMf�TK1"�M&6O��L��J��ˠ����Q�x�-��k��!�ȿ��B͜x��GB� ߬M��E;���zo}�Je�:�t�\���c�yd�w�!Nȓr�g*�LWF���T���I��z����{@���4��탲��W67٫Q
��9fn'&�������"�h���MxN��@�d��jx�g~#���t�9�Q��%�3�)<�S��:,^+���9u��vv�3|4�+)>9:b-ݱ:�}��rF���zSWD�2 ]�X�a�e�UM�z���ʘm�k�k��_�����^�dT�3��@�T��C]'=�]]JP�ه�7ҏ�.8��>�ϭ#y8���q�x*Ȼ)�� :�S�t�V�9(�X!��j>���� zi������}�a���NxB�R��@��@�� ���m��6a�}dq�L��wܪ�@u�wN޲�}z�ܢ|:�w�i�e �=�'m��#w���:�4DI�e���hG�����r��\����{���{P�]�\&�oB=�w�/O��;�+�ھy���^�?�f(�t�B$�1x|d�H��+�;Unu�E��#_�W}�����]��s�R试ﾽ�Y�kRp��x������}�dѧA�����I/y�q�D�Myƌb������]��3Q ߍr�>�Ev@[i��R����A�I���9�hW��6�	L/�l���5c�D#���U>�LēN��[�F(%���?������8����4�5���xWt-�l�&N�0�:�q�7�҉���wE�>�;��*)V
 ��mdZx8=[��d��T��l!@�9��d��n���b�L�n\����j�c}�h�i7�p�Th��p�W4'!S�����F�8^�)`UO�o�-�w�5o�������y)��>���K�������)�z )�ޏ��L�r�<����ˠ��I�}.�� !; ��a�D!��\w�������[�Ŷ�������I~�\�z�ܻ{�ܿ�ܾ}�[�L��U��Jy���+>����>H��u��b#Z'��ӣ�4\!�?٠���F�jw�Q�u�GnM'bH�!Є�@���O�c�O�����9����l?�S��X�����K������Tz�}��42|:a�8��q��48A��J�.��0]���A߼h`�t*���>8~��5*�q%4�&nU+��u@nPp��pp���AA��G�z��߶���w�Nݻw�|/���w5�sZ#�u������uT�-m�g/ޕ�B.��9U�P�S������� �/��j����e�[/�;>(Ǉ,G8(ӓ���y����]�y�Rr&��ػm�e)�++�ʃ���:[D)y@���׍�!з�
�n���r;k�A`�N���}�y��@I̼".�ڻ�4����)��a��Ŧ���4���)����Ն�t�!v�SyK>�c9��M���g�"dA'�I����`�P}�h��\6U��_��r�'�[67����Jy�f�,-��"y6Ecsfj\O���������I�H���`O�㞕;*"OY �������@5G<0�*���V>�cK����0�u+�7��|4/[�-.m�#���b���섏`�����7w�)��3�<�-���j��h��6��8VE�.>0ʅ#gky�g��ϵg6W����g 0��_ �_T���G��8D��zя!_�t�DI�z���@?H�m�S��"��g}�Cg�;B�|T9+63E�:`�N`�Оn� ��>`t�u�|�ʇI�_��?���6�6����Կ�)�{�27U�����[�����wߕ�wo���g�����,.�I�]+���)/^��N���>��ê�4�2����� r�qܢ��S�Pn��b����8?]�ܺ^~������^,|Oq�K�^�Y�.	�7��6K�b��h������,� ����~T�m)�S��-�N:rw��m�ۤѱ��.���AF�{f���u $h�Ƞ2s���0��%��q}=��Z0;�3��M`O�τHZ-��� �/M��crGѴ���r��"���}��{�#w߼],KK+ew�-a�+��رpy��oo޼$���'�J�p�Ӯ���<����'q���@Q��X�!���+	�);�	��AỾ�㓼^�R�[/��� WtB��r��e=�����׮JɟW���ၗǼ?"M彷׉|<&�<	��k��Sg&�9�ڊ��>�  ��IDATj'e=H���?Vn�����{*vҋ{g���j��l[����u�mB4�N�%���p��ُ��?^2�� g:��݊-�*= ]��j�O��C#mY�y*o5zd�n�������G,}��UpNB���m�#����Y+v�տ�S�})��e��x�����o�￻_�ܼV.�s��Xa7�ͭC�;�������E��7
L��)�������|�Ą��s�	�Wvk)�_���
�p�f'5�]�2�ܿs�ܼvE}��b��B���[^<_*Ϟ16n�{�Y��I���[�	�wώ��"�߇_Р>5Xi&]ꝳs@^W���F�������Z(ŀ��Q8Q���T�^�M�d�/6�
�+�� ѓq ��t�����Ur�/[���c�]Z:��9m�wBX^Y-/^�z��O�9�?r��������]�-��\-�n.�f.ϽWvO�-)�jH0A�d�t�1:��S�@}d	:H�4���x�EQ�g{s�������u��ek�/�?�:�N�/W���^+�>��|�V�]�P������P��-]b�n9i�]˄+�zE�������Mܼo��3��V���ʠ�~� <3c{��L�L���t>�_�gM�B����|��B�Uo�J�	S��`m<I�G��ͧĆV�/�J����䛁>|�3B��q%gR=L'숟N(pP���n*�n˲3Xq&OX� ���?(�S����r��B������wo�|wA�����9.���_������������r����+�r;?2"�Í��'q�_�n1c�es}�?e�>��EJ�ܔ�����{»����e~f��)�Xg��vX޼�,��)Ϟ�.�Rn�vE�}�cI��V��RlH��2����04�j�?̧ ��s�u�m;�)�����ok����@Zx%���L3�U��X�^�u�͊��f�Gb�ۭ�}즼R��	C�8JE�kz�Nq��$ȴf~[�,��j
,�U��C/!��뤼s��Gꬶ���ʫ�o��nmE�E�859⵷���e�/�y�5G��HQ�Q����Ԥ�y:8����.�	�M" z�?j-�Y����J�z�f�ãse}�'�w�:1�o\]a�1O�l��'��1u~��^��{K��r�´:Bu�R�5`�F'�?	Fz���ν/��V`�Y���(��psG6���������G �A�?;�8m���Ɂ�@��o�W������N�����f^�'U��́�ۃ�Q7�4����M�s����m9�B���s���`*�⦥C��,�(�}�B�/"iht�'���O�ģ2Vgl�ӛ�����vv�ᕼ�%�������/o�ؾ,/^,z)��ŉk�N�J;�W�l��֟E�a�? N&Hޚ����<��GG?���妔��%����g�[B��4&�,oy,x�r��{����� 0@Ͽڪ�����ٻ؁�R*#���� y��u���J-̜����:>mo�p3��QGm�[M:�HQ�6еN�*��Ci�H��q�6n�T�%od����D�6o��a��^M�Ri����$*��`�\��S��Q�z�ᶆ��2뢤`�K���Q��ZEHG���_�V��7�����*[��BE	��M<�Qnܼ���	�])�,c�U�j�Vp���*t9f���i��{�?���b%R�`@SW�<���4�L�T�Ѳ�u�u����*Ϟ�)oް��@�?qb�sc�֍���������+W��NN�/���;l� ���C�Q=�,D��V!�I��F��2����ӽ"�@�ԇ����L�c�FN-�l�_+1��ap��� >��<v��F�ՠ���	��'��@V|�ןzX�v��|��h��Ue��9X��0o2��x�R�.�m��h������ ;ybE���n|��X��ۓC��r���7GV�D�H��a[f(mA<pX�y/��w�Z����w��)W.��I��s�He���v���_{g�'�_�����^rL�Ζə�261a%$���j���V��_�iVl���$��X���B��ڮ~��?�u몷<�~����z}��xǷRl��m
o9� [�C�E�*��*����3����u#�G��š �a(h�`����qE�hs���t�<.;�t�_����:���j��pm��!���مa���7����n��Ȉ@�������|+$s0-x�٭\<�Q�N�N�{�Ƈ	�������O@:)���*T��M"AjФoy*ߍ��u#
;�C���M�?1\���	߄k��{%cm��iĩ�W�6v�a���'kO��o�w�k嵔�wKk>���W01>Z.׵�wn-�k����$��Q��J���-=����\��p��YpF��[)��<n)[>��c��Q���5��W�_޽e���^���n�lm�e���+�c#e�¤��>|p�|��O�aV���C$;�ȌuW��m3{sE��qgB	58��4jZ}G�>߾0�;��ܚ�S�){��Ue��ǯ�O�ύ7R�OEAֽ>h��p���2�`t���)�w��?�?��_:X�rrY���.�@���?1K�`R�{`PЮ�7�*va�� �y5��v ��r|e�
-�cY��^�v��_Ԛ���2f��/m�U��h�X۳!�2�x(��}��oŀu�R���h�\�|q�ܿw��l�yp�ܹy�\���.9��N:�K[������y셾�n2��Oi��A�-��N�� Ϭxx쯼Wތ	��]�#O>z���شկ���P����%tR���|�ܹ}�ܓb�vgf9�r�yƒ�������jy�r��.oz�[�/��I�&�v�Z����SV1\'��=G���H��X��_��j"������\�G�����W��M�rY�����Ӊ��V��R� F�ݦR�!��@�`�wluY��\n��CE��rvp���뿡4�p���7ZX&W[��%Sc��X�	��i��^p���!�q \����5�V��L�yDʇO)�q�Dx��m櫣�2�e��5x	�O��4`>Уa#�e�)׿�!�Fu�7�=_*�� �H���<P؆�Zd5��l� >E^��$�;���V�M�FGO��c	y-595U.^�Xf��U)x�_b����3���]Y[-�z������h���+%e���7Y�?�[��c���bw�
U�D_I�	�n�A���(Uo�;����N+��&��'��6��UF�cc㎳��Svwv��^�b�rʛd��(J�NVi����.B��x]�b�;/Pp5��ty�&d���:B�k��)>Ҍ�D���M$���u�:� �� 4D�c~6����O��z�ϧ�h5C>�(�n�� a��g��$5��C��V��ПKQt��= �]o�T�cP$/�0c ����D�@9d�} �y���Wx�[?TZ+X&�.�\�2ǣ@�0���9�������W��e�poڳ�e��2��w�墿!,�䘵���,�����ݫ��ӏ��{X�߾.ewև�
���N����y��^�E)x���B�<c��>
�je~�)�Ñ���ǯڛ�^ +��<�y� ����A�r���֕��R�}�I��o�������+�����x����C���P^<[/��ߟ�_}�[�zv��2�������^��ܻ� ��`�cb�\�ކf�\˽C�����RL>I�1\y�@�ژ�Ǭw����h�Θ�I���+f���8����ޥC�N��IO��N��	�t�C�D=��pϏ"�*[��gtѹ�G��m¨��PdA��|[�{H/lk*�>���Pv��\�r�b(����#�u�SL3��&���R���d�L	ɤ jĈ[[Of�_�pozLY�� R��E�(�}�`A��(�����'ЎG�S��(��KT�_�[�}P��bT�}��@Fn��_1ﳓ~���-8Wl5D<��tt����Q<
�-+7��z��;1>^fgg��M��#/�8xM�{Rp767����Hy�����E��]YaA<�l�1�jo�p��i�1)M��vL���� ���_��cW��ݕ�ǖ��xQlQf�x�7cj ܳ��vw�������Y�|��D; �	����.5/���������~-�V�BڻnߊhǙxM'a�h�y߅�qO�Kl�� &����pF�=y{j.}&D�FR�X�ǁ���I�
�u���%(����`��Y1�_d���(���p��Y2\EӨ���
��U���@�H��}�]�������3�s
t��f?d���A]<�� �/�W�G��Ѻ�9)�sRl��^(�}wW��7�Ὓ�r��e�d�ovx�b��������o��7+ekk_�5�2��0n(�Ш�C���P͞������y�b@�����,;}�x$��t&X^����y��)�wʏ?<,wn]+�|D�>����ny�h���OˋK^�����x��~�3o�M;�gH�zƾ�m�׹��$Lx���p�l1�2�t�I��~sW9 4��Bz�u7�9��P�G��vp�"1^�U��������1cZq�c�'��/1�E�%Ѱ���$�.t�x�JVh�̎M�����26)׊��Le�������[��-&G��z��h_c~(�q�������b#���h0IE�5����I�"�T\Q-T4�"�ѹL�@;���D�U&Y�e�V-�Un��.�\V ���b�WA��� $4����y)2�T-��Nw�Pp6������@��m�n-f:mE&L�c� �[a�f�І�NN�0�c�6~�A�<�df�J�W��Rrq;>�P9�K����7����'|7�7=�NZ�z����[fA�<I2�Ia�m;���7X�I��� �vt�+�C�bv�Vg�f�@џ��Ӡ�3'1Cqy����*{��: ��軆!��)R�qR��<:b#�c�+�;��͟��;V�.�)2!�-�.��W���>2O�
�τ3�${��>�����4�����,�O��E�T%�Ql?�Dӂ��t���h���ӹ7ϭ����(�4ڰ���xsDC������������s�/� ��D��/ɎR}7o���֚��]��������� ��~�w�F��A|J
}'1���_~}W~��My��/V��ڎ?:v�%ެؑ�0��;��y㫊�/N���o�n|�@��˲f`�쟁ds8x��H�Զ�}���~}�|��})���3t(:�w���=z[~��Uy򘏫7=��~3*ō���f��������h�k�hE34Iw�{�����>_��7�]块	Pg��S���5�x�ӊ:M�7t�(�ZVpG�+1�3.�rjjڧ����[sE��c?R]��QnAٝ�.��яIE��,�2�
�t�����d�
���d��&})���v���Rz'��䴔_N%=�L.��`Ou�?���0_�]�r��r��*�Cf�95�Ba��!�1�R$�&��cj6��_����7W/�I
�]��j�J'd�:�ĳRKg��ew��/e��&�*��o���@�^�������@ƴ�1]d��䯛�)>�G�*���h�0���Z��I��dR����'�}�v-E�`{��������:���NB����"Ws�0�h�ސ[�b��x��^f�y�A����v)�4�=5�#ֶр��9�L�_���-��ӵ�����H�-P�+�ob�<ڬ�m���>���I������!��J�>�H��4��>�K����7��3!K�!#�^�S/?2>�����Ύ��cOr�z\Q�h��צ;�fߢ�.�/H�G�p�I?�F��'~��F�����1W}��V��>_ny����ۇ^g{U�7��5�x\V�������y^~��uym�v���J�P��m(C�e$/��.��r���#N��{d<����f�;�����7�GG���T�}�Z���o������\j�g�fg���~�V�"���ey�fų��|H�D����| !�n��7��f��5� �eI ଂ=�Keh�Sz��!O.R�1�x�7"@�zVu#�F ǰԵR�E�� e�,����O4PhQl�<Bɍ�
�б�V�b��,0��.w(�{��[D^�	e6a�	F+�<�U)Gъ��l��2>ܵZ^(W/_,�.I�����߼��%���������%DT�V�m��ߢr�f�����m��B��-��X���H�V`9M��ɐ?�H>d�q_)F:m|���r�{۩��5Z�PP���Jw��k,)uen��\��֓и*�z*��q�+���Q6�v�RYX�#��KT�d�8$TÄ�@����W�j�K���`�KE�5w��sfU�����K=c&֯>h�n,Eko��f	J���m�q�@�|\F�n��Y�A?�.�<pJ�{ӱ���y�𪀧c~�P~梦�<���σ3�>C�3E<L�K�|Y����tp9����%���� ��'�w��Dv4��|��u=ӤJm"a3|7��^C��j���p�IOfg\@��zB�wy���6�v4`����~|P~������I��#Y�oY��+�>Y,��y���<*O�������J��J%pi�C�5����m�/l�����U7�FH8�-aG7BD~e��1+6
��jv�mz��ƍ�偔��X�ܾ^�y#��=}�����vy��]��??�����l����r~�W�R�D7��`�\�4vܒ/��#`�@�[���{�`ܡ��נ#U]+1G�v�Ue��Q�k h��U:�V$��Z7�|���Z�A&�x۫�q�rk=K�"���<y���G���*�P�?,=@t��e��h=HQW��E��VwES�� �6Œ~F�����7A��mG����b��N*��1�w������l��2B��
l:�t���e	.<ŏ΢E!R�\X���fE��"�S�V�q�7Q�_{|j��#b�pK�.������Q͆�xg[�(o�Xr�g.e��8'|m��힔�C=�M�ʀr������W��Mv�Giј]0���8�t]/E��<��z�W]c��$����S"�sX�Lg�ɒ���T���B�PJ��#��-OXy�p;ѕ3�Qm���W�o����ی��N���)^@���A��	�p�@�2��>L�K�|Y��u�Ӏ�_D�u�mK)w?~"�|'�	Y��^>#\zF[��՗q����	��G�axp^&[���'pi�� �nd��̌��W��7o�?��[���8q���k��9,�����e��ߞ�G�_�ťu�_RLԟ o��(��ry�f;6+sM��a���F�^y����%����Eh#��D_���R~vg�\�4m���o��(u�i�k�g�v�Y��+��_�}R^�^�΍j̛�GJ(n΃�V�.Z1�/��An_(/��s���@�a�HRv`�K�K?r7'�����PT�t׺�g~��B�c,�6t3Ygk���[OjV�`�����W�0~�W9A��(��̭�?dt�XW�'��~˃<p��2��U��,���q��\A��r�)���i��f�D'Ô`��5K��!��L��b(;��в�δ/Qn��$(Od8��A���t�װv��]�ĭm��W��P��?B����4��-]�T#��J��)?��h����N5<0S	p�p�W׼s�Ӏ��Haq�<�vN��7�oO@���]H̮g�w�}t�8��3K�u�*���ݲ����05=S�Y[wQ���O�/�C�e�����A��R��� (R�p�U��&2O��!�G���yȿ*��^��@p�S��z���	g�}����`_B���Z���"
VN�>~
��������h'�����7�����c`s9���HSP���S�8���g���@�˟�o��~pW��'���p����ߖ���a�{���q>��~kۊ�V��ѻ��<�b��,�[�b�>�5�<�kL����רs�=v��Yi�	�}�Ha5���>w�<�C��r1�O:F�M#v�W��ٹ�r[r��wߖ��޻%��´�y����P޼�,��y��OϚYk>��#2�p���d�e��"]�K����e�J3�����%L]&Ɲp#\hU��Vr5�-(�L�����I0�[_�	b�t�	GPώ���2
CQ��:Rp��<� ���B�S��֦b�~Ї� �-�BCK�E���)�Q��w3�{����8�ہܬ�q�Xy��K�eVn�_�-��۲��L�����F	r��A��_UJ��rb:C*=ϸ���ܪb?����k��ԅ�f����3���<ͫ2�G�%�S2	�
��Q2��Vle������ZQqs�.�������i��yox�5�I�6RB�7���>L.��Y�'0*��
~_
���R�X�0��	^�`喏̤ �3\]]Qg�]T8Ho��|O���1͂�*`������pk��� �ГE��,��s�x��P�>�`�L�!��S�|p�,
k����+/��'B�Qa(�r���u[1#Ȋ_��<���~�0qA��F������j��L�I�#������ϐ�ĭm��r�"��d+�O כ�g�Y��_�=��S��T)�����Od�D;!j%kg̊���#�c���~	�_!o;NC�����.f*��g��1>��xi>*/���c˩���ʔ��\�P�߿Q���o����!<��ŷ( ��}��Y~y�X���+�/��7+eg��[�,��C�gma^H��(q����O��!���`h��<�'�!�y	���q�XJ�N��Y/cʍ��}��ܲ�¥�299�{��eye�<{�\~�b���͗�5���ϖR|�T� sr� 2������t��}� �<�dE>��	��ƺQ�'��1ʨ��i���y-3��Ah��S)�P%Fޤ2k��
�4A~�����v����=�����X�K�`�;�e&%�S�y���,1[[�X��h�I�#)��V@&5�6`RnET���n	��7r�ORn-w|5��f��'��
�	�[h��e�G���ؾ�D2��L7ˢ0�F�ʨ��;��;�Y�$�p���c8{��"��R4Q�� !*oA�Y`��)���$7�&��?:�4=�Y;��?�Ww�V�/�l/Ҍ�͐@��;��_߅�6d2z0!��KaS�&�ʱ�'���5(55;U���ʜ
zZ_��'��ĭ����܉'#=a�<q�U@�^�"]�X-3F��ڣ5�q���fK����V�t��ίIŸ�s4 �((��ƃ9�לc���2֮AN�ǖ1����%�����W�=
t�Mr�딭���u���w�h�g|;����c��'�4	�Ѿ�@N��x#����O�A�'� �����4� p*��G�'��NSVԟ3�	ۉk9d�Έ{s�H�4�|�Y�7\ɇ��a��Wh�c6��y�>����q�0�S�-V��V3r���4{����8(�}�Jڞ|�cQ��Y翿��yO}��r��L��������;���9>��XF?��sX�.n�G���}R~��ey�v�lm�V����y�ԑ�yG��bȕ~&�ͱn��һ�{|�JT�M��#����m�0��^J�����bK��[.]�.?H��K�g�捅291fz����~y�l�;$����`Uc���������&ώ���#�l�^����M���y���ş���Gu��<��Z�Tl��"C"��m�9�F�G��1f���C�-t���_(��tZ�5�����k>T;�;�@<&"���-�_�u�����z���)�lvNuf�Yw;r�(�
��C�?2ӷHo�J	ʤJ 1��^�y�TB�L�i� �E`Z��d�Qe��Mdܞ��N�m�EHţ�zfn�G����6�T�( !2�Xy�J�|U��>�ai���&\�(5��@[�(�ֿ���{E7��#m?d(���ٔ��23;]f�f�%=���L�Q�<P���nK�E��>�.�����f!�$י&fã�NC`�;��Zh������E��\k8/2y!�`8��^��en�#����Ff�ň�P;�)�JGCV��).KBհf?y�Mֳ~�S�7�E���6�_���u��`��"�4y�y��C�������@ PӠ��EKp8���4�붴>��ׁ�|���� Â;X� x�����=ݪ�gv�u��댼hH��dQY�P��u�Nr�X���7�ġ��F����:fl�ݹV��BQ=�>��������R���W�??+/_,���]���ٌt��t�0cd�}���(��#d�끾��|B�A):5�!�ܭ �C�&t �=���+�S�˭[�����=�p�3�,�<:|_v�˛7嗟_�_}�vה/G�eΝgbk��4�D��F�,�eInݥa��3#б��� �ҟ���`%�<���x@q	]#D�#:�|R��Խ�D+�<�.��ʑ&tL�t3ܬ\
]~5��A����k�����	�����RnͲT٭�V��R:�m2��6�D��˺]ђ�;9���9)��,�����Pn��:"�4]K ��-�� LdP ��0����LS���-�B����fP�I�I��.�3e��G��`�6��,��aʭ�p�jx�B̴������p��|2ؿ���jW�q��i�0{1|�J�ܪB���ʨ*ߔ��gf���K�����%�̍r*I*�;{eW
.v��L�Jep�y؈��"eh`Ի*O�	:�pD����O�宗��R�>��C�~�qF}��,
���[>>2;�Nt�'�MN��_uQy711]���O�:�b����]R$��t�;v��&?,�u8�	&u��B�˼����D~�����@�Z�O��u��~~�_=�"��@M��]�,8+���ꥱ����&�������	2,x���G;
ɻ��>��G�=3p mQ?n�0������ّ$i����9@ �IfUvV���,�ڝ��ݽ�}��ݒ�ϰ���$���; ��~�'"fz�w� ��]r��2QQQQ&�ƀ��~ίu�����=.�ro!���B�ƈp+�������s2��[��eNSW�{�i�FF��]k|n��ç��s�ٙ|7R�.2�y�,�� 頄O=D�sE9(*HfC����:<���V|�"ɶ�����I[�v������O��܎���r^�s}�ߎ��?^i���<\���x�>���;z@��^\�$�?�.�0K �R�PNRτ� yk�A�]�6ـ�FN�Dӿ��򚧟�m{���
�k}�6�Ìl�oս {��b��!��l!��tH�%�F��ʪ���<$6m�Z�e#<��ed�V���''Z�5m�m	6n����m� (2�91|&*X�d:ϯ��A�$����)���:-�+��{���1Yq�����^��۶&3ފp�ރv���v�>l�}1�[n�.�n�|z�}x�v��ɶr���L����\��q��D�g���N`2$��i���o��CT��D&��?��[P�k|�����Zn��z�������G��S��d��C�g����n�ϟn'O�}^�00 k�v�}ګ�L�{V0 �˛�~n���/�&���O����E{���lAJ����;sxІ� Z�1y��qW�0o����8x@�._���}����϶�2v��,Y�9��v_Fܭ[�ڵ��4�?hO�<�����m��j���G�P"��z3"��~��U���A�@�Y�	�
�@����@�0R�o����̙c����ٓ6X�D��mˈ�����yܮ]�ۮ^��nK�V׼��4ϳ�aPizv�����!��2�����H��+��ψH
Zߢ��.�N����X��Pe�S�)���+���h$�I��õX�F6^A��h���ax���o!� Q�C�U�\Ѝ
D��AD����-�eK̸NU������ă��C"n7P+M��q&nP�Q<��V<���Єp�A����v�ƍ���K��lV۹sGۧ��k_~�������G���?.�q7gZ�9�U��y���!LWHy]��'���	�5!�IBf5Bq�,�*Yn���ڽ{O�?�ҙ���/��n�x�?��m|�a_;x@F�ѥv�����z�N���m��QĘ&A�����R�n����o��?��8��@�E@�� L'垝�g����{�p�<�r	P�}�����H�7|���v��J;���W|������v����q�u�<k\����.ޚ�AMR*�ڌ��}2<
˜��K����`��0t����)�`�I�2@�ljskƑ#��������f��8�NKk�/_�'��ڭ��ۍ�wڝ���N��5N&�qA~w/ud���:�N��$��AN��%Ht�-#~����H	��i��{[�p9`�����5>�DP ���t	���}�����%����@İ���JSyv�e����> א���9�Do�i9~�\P2u0F�d&n���B��%�,�\����rڋ�:��Dg�7�7��{���2Z��mn^1s�����'��G��AwXͼ9�T"O'bԩ#�Y�Y�a�dL������Sٵ`D�tod����B�eMf��&��Z._�����V�v������ńW�,-ϵW��ʊ������:!A��a�3DL��K�?+��7�π������S�U}�?�)|������,agl�Y�o@X�5�3����w�B�!]X���؎;�Μ9%����m��q�k�\mz���A�����7۝����*�٧��{le�b@g�)ͻrb�]�4�)ֻ�rY����rx�� i����[y�d����\�o�Ȩ�t�?/|�S��nGඌ��=�ѣ����G2���2lWW_���s~�dpV�s���^Az��-��������ժ��y�_���p�:��ҷ�ض������q��kR�X� D�Ig�%_��H}�FZ��;�.�T���@Ũ���0��t�؝��:s�$��I��!5����:��EM��)��"���?(}/~L(=�A/�,,�=o�cFT=x���E/��/41����x�]��{�./��I~��,�/�l]:�	�P;��CW&ٲ_���Q�"dy�:�T�(ݼ5@Z�v��@�Ǝ	X|=��/z'{a�@�?���7Z�u��+�����?���W۳���S��}�0e���o\�$����o���@iN�i�8�U,V�#�P���5�=���a�?w��S��`�(�=6ӝ�_�_f��M�1,m`���*ɕ�c5q����!˞0��aiU�\�1
|u�)��1�8v\��Wڱ'������O�Wß��[�}�|�]�q�}��5��s�i|�kcÐ�:��mĲ���'�7���}���G}0�皎����W:��ޣ�zݔ���sí 6lU�}|<h�>��+���w_�/>���?w�o��\���Ǜ���Wn	�~�$����ۊpqyI|�Y�O��:�:���~��u��<J:����X�}j��D ��\�Z�@⓴�=`3�������"�q�t6��[o^1\?�s��S�(L���k���J��U^�ؠ��u�b�\n���z�-[$�[pp�>��
��Љ��0Q/�Xܝ�������2<�`�i 6�[��>��*�I��ĥ7d�;��R32�lFMP�K�����c	̦�S,�JM]��BX�ǀϴ���`���60;��4�l�N_/�̷��������vp���}��{�ԩe�./̷�GW����ڥO�k8Gu漴�	�>;
��X�� =�t{QPY�|'�`�.E/����}6�B^m�Ğ���Y�|/�������/�]o�]��._{Ԯ�x�n�y�<z�Vub��Z�������C�(�e�$T����+��v�ͤ���,,��?��J�a`2�0�,�56��w�ނ�M��]`����*j�Y�x�g!�PF��!iw��ރe��Q��p��cHS}z��N�&������p��4Fi���p����C�4�i�E��x�u�E�I�ys{���A���1���P~n!�؊�'�Z'ѯ����Ls��'����U�M�|u�/�\m׮�i<��S�����ט�'�]+�$���:P|H�߸v�q!k�c<3 ��a엱�Ʀ�(��Z�,���R�2b������O��|���_���Ϟo��^�+�﷫7�{�z�F_|V~���+5��)�D��D�)���OYH�1bT5�f6�N&�Ȓ~XN 帠 �;��b��|~����Uݪmis�	}�-Y0���� (,e�w��7,M2@�/r��ڲ̔�O�*�dHZ\�2C&�v��W��J]��<�2a'\�m4�qEGP�6w�7��?X()i����T1�fy�AĶ�P7m�)WB�B�����o7 %��<`-W���>\5�Q@g��(�� ���!CC��~�8R�GAY���`�c���T�v�|��~yB2_�%o��p�7E��u�5Ij�q�\���a�IЗ�<H�8�V��ۊ&>I�{�ԣ�v|��ev0�_���� &S�:�8�!,�Q���g¨�ECFD-DC�~���+I�q�D�p!4Dz�\^�����Sj���[[����ɶ�0O�o�{�_��?7o=iw�=i�4�&M��K���ȍ�|��}��Y �\�' �d��ŀ�<����?�`��q��rVz������c�lP�҂J�7�>�C��Ĥ}#�vG\�{"?��Pr��۠2�i�w*k���-��ӝ<S8ى��)��p�t0a�]�J�Χ�b:>��f2Y����H�XWH
e&F\���?q��Bm���w� �;���5��������8��R0��r��r;x�P;r�P;s�H�_ZjO��������[���J����������Z�T%=֮�8��a��D��gL'T,?d��x���{��'̒�[(k!)K�#�3Ӣ�m�e��}������/�������O.�SǸrȃ������k2��?��kw��gk��_e=��J��wl=��JS��{�}�c-�uSs6��I�V���K4������q&��J���6�ٍǦa�v�Yg�J��*d}''���\i�U�B�se��`�v�]}C>�1l6��u��g�\��,d�qX����IP6����`r�f],��!_�A�}��h��;��]�Ͷ\oK8�'x���s_�_� I��̌<AD �[*�4�M�<�Fd�Qt,"Fc&_+�7n5lܪ�����:&��Q x���BF&��-�]|x	#�$���Y�p�U`$B�D��M@�ORP7tը#���7FC ?ǹ�E��!��r�Ty\����$�=��!|jk����W�ۡ�~hJ�#�/�P�m.�3���/	��B؆m~`�e����Ǯ�c�?i�ʡ�;��v:X�~x��!N�!�\E:A�4��&�M{m|�l�=x����ǰ}���vm���Qy|[�u!Sɝ���6 ��F�3�|���d��C��&ܝ����G�����4�<f�#�fa���:솳3�(���	I��7Lz�����a����׉<���w<%�w��L�u(��>�9M1�c���t��M�����$b����*lz��g�`=�TD���& Nf!F�K�Ҳ�f�Yr	/.,�����mQ������굇~����ߐa˭Oe���n����Z���4U.ŀ�"-0#Pd���-w�<F��C��%;r����b�����K�k
o�����ԩ��S>Z��G��.�sgN�S���2�<^oW�>n��p��߹���m�j^���2qٚ�@a�n�������� oT`
�R�c�H3�u���.^�I(;�E�*Nz#�.��I�618�AU���l�GPB�3�H������H,���l�a,�`���!LJ�C\���dڀ��b���e�<٧��������ANҩ_|����#�y��6w^�-��<e2'wA*$\	"�H1�9���"�8�3����10D�l)��-�,�'e d2Hީ(J/��2��߄<@�Kh^Ȇ?� gF�̤@t����,wT>�DmG_�z"$���;@ny")�	�YŤq>�j���O\#�$ՓO١��e�\�܎�岕���w*.�=���<oؿ`#��<����ܒ�1�����;��Q���qC�{P���w�-9	�Fyx�ӥ�GƂ�+�,���@�9�E�/���ǫ�у���������U�`����]X��y�S�h[ߗ������!������<)�@P0.� �OƼ-��a���mT�]z���I��$��+C��̀���| _���aZ�Ӭv�i�.��g5Λ��;�AU�:;��,U���"gڌ�h���Q���ư׬�X���I���i���
�F��^n��ɴIO<BqE��0<z��ݼ��]���]�qO��:�~Ԟh�|~>��U�u��ѡ�cQ0oEd�1���Br<�7���G�w��~7����d��y�𥌑}~+�ǟ�o_�q�������k�/��^m����q����t���,��
r�v?��'���NS�a?䜊;VT ��b�Ϸ�U^a��
S�U������!���Ua�4�2BՕ��m�$��.�[�e�n����x����n��$q�o�p�T���<�t������G#�E�ߴ��eܺ���QhY�]!��#�ꤳ�_���|�>� .!�`����`����wv+g:H�����Q�N�$\���!�8´ @q�D橊8:��`
"A:c^A�H�I�ًv��v���v�W��yܞ<}�I��'����Ξ>�>��\��~������7��$֖O�//��c�����Ff���>�w��q����0���f� ���`*��y`���^�_q�F{��y{�����'���g��sޡ��C�H�.6y&���Ƿ���}�{�e��eE:ę�ہ�I{$�����E����ת�t��Lw�i�	��-�=����И.W��:b5�<F��P��S�#��C�3xN� g�������[�0 �?���}�~��f�˟��ﾻ֮^�����62���� �v�ܱM����,eL#���>=�'d=�HØf3 ,Yy��k����v��r;�T����P��b����=�x�͋v��C�\_�~�=z��ֹ=L�c���[~#2��] t�^A�j}��W��D_���iF2\�hc���-��3"���7���a:<ނ��=ʟ �wZ���ۂ�^�����w�j�YP��� �8fѓ�	����qpq�
FO��l<��3���Y�&���6��U�C�۹s����h}|�}p�x;p�]�İb8c��-�yv4� H�6@���\
"�+ ��c,}N�0O�'b;��h<i���u�L6�u&���l�{j��]م�%��}���h�.>��f�RL�}#P��t��a��l�aG\��Ll�P�zsp/,����:�E��؅��?D]ug�w�E7 <@ÿ��@ԮbU|�>��;A�W{���c<�Ƌ��������C�X?������%��ڎ�iiѯ$�WZ��<�Y��ل{�Ҧ�v��i��k��n<ǀi!d'Ԩ�R��m�-�hgNk]�x�����۩|�v�o���nܼ�~�Ẍ�ۍk7���Uo� �-���c1\��]v�^?'��[��u�֞���.��c;�fM�P�,PժF��$�������^�/�0��q�7�h�	w���xV�qY	a�?�#F�ȗ�-��b/_n���q�~�N�|�F�r�v���߉��wx��b;}�p�x�L�t���ڱc��Ƅ���.�� �#YB�< ��z���2����#@��"S��;&��v&�YX���C(v��]�w���0�O�ÂJ�k��<ߧϢ+���~5p�*�o#�\�Jc�s����T�6�E��=�A���lCŌ�m��Z[_[kkk/m���M����
�QL���]�`��{�a�c�{��$�w!C�zů0��r�e8JP����}��A>�p�]������sg��cGڡ�%����O����w�xM�r�f�s�~{�a��W��9o��̳ �]����u(ք:�����h�q.'�7�u���?�]3��a����¤�O�Ÿ}�0�?�"b+��ΰSX�ηG�#i�r��+9]�~{|v��vy����ym�޻���x�z���k�H��9y��,��O�/>�Ծ�������ƭ	���-M�[ܓ��;�~�+4V�b'�4F�(�{�wx����7`�A��p	{6�Pi�c�Ef���UO>C-b/4u�yP���z��������)��a���ً���/�p71��p�_�4���^�t�_�՜�����Ӌ�g�
���}+�h]��\o�:8s�é�qp�g:,���<3�}�杤~��0hƓ��;Щo�h&�N��S�!_��`�V6֋��y?���'ZK���}|�B;s�x[Y�_�����n�y�~��v�����ƍ�m���8����W|e�:�L�{����w+���-,�<�{��[���`ؖ�8Q�5�	G���gl��Sճ����t�+T:�c��$�8`��Ƹ�:�sx�L'������ţ h�j��Cx��'�	0���184DMeR\%!�ILi�i��xP�Bh+XЅ�,J��&ژ')�|�T�M<+m��~M��>��k�d��i7n=h���h/��X]\҄t�?���z��уmq��D��!��0�F�B�
G(����,�$bTN����A_�ku9���������)߀D�l����Ã�M����r�w2�X0]?��?R}|/��U�X�;�+0��Ӳ��3��_��O�`g�A�ෛ����;�-���9*|����@���=����F��r����K�}K���e��}B�� �����eɿ+SO��;串�6�!D��31*�hL�G���d����t;t��!������x�onw�n�.��2fٵ�t����ჾJȴ���=y���ڕ+w��wۃ�O��ƶxq;ؼt5���FI�o��$ NB��Y�����_,홨��-Mh���CEȓc�x�8��OA&'�NpY1/�ePVphd̠��	��� Hz�ސ��.���?P��jU���H�I#tǦ��˶s�s�{�L�u �a~�'x��'c����3S^����Q|(�?��\�����H̋3X��s�rՓ|Bn78�0y(��&�|[BJ��(w�RDd:�H#*;���G��?�i���N$w��x�h��Ge�<ЃxV�m�%�|_�����hd�..h���'!��/��3$�������������v�P���QK|R��I���萀6P� 7m�h�4lE�ab����*ٺ�b1�;��«d����t^�,%����� p�8�ʛ�<����
J�A�,o����IL&�Q����`�G�d���C�[�c|Ry��x�H8��B���Mt�o����i �07�T��̿{��`����7�ƈ� ����b<v�y>���><ƹ�C��i�/�Y�.i�W� ��c�@q�6�qK��p�1��̀���n%�f��+�,1��؎�C�ɼX�����u����O����O���Q��BA� �X���M�NeMb��W��M��덏5�v�3g���.�k_|�Q����v�o�Y�n"��:��[���
^�v��=�5/�ƈ�_o[_�<�Q�6�F��#Wul�pIj�����C@�	S������l�k���b�or�ITS���'��#��|&@�>Zn
�n��!?�cɉ�����*�SV���v�g��:*�"+�7�,� u+$"�G� x�sI�ޔoK�U`�#>���mR�	!�;����_��Y`1�r"��[��Ec���'_�;���~w��8`��g���i@ԡ� 3�I����0� @]^��}��14
',{���_�3�ȍ�wۏ�niR���?x�^�����e�>��Μ>�><B�)����e��e[��&}r�Q2�.i�FT�/����ȇ+��@O�aLhcZ�;��W�'��#�F>1��0��6���'y⌼{4��:M��`/��=aB�]a*��%~'o������v�`��=� L�]@-��Y0#m�_Pp� bd���"2%�!�v ��i+n
*i*Y%�H�!�"�Ȱ!=D:Ms�	v�*o`��Mؗ��6��2�`k�͸IO�ҳw��u���.��+A�X�*c8��ج�i�����3�4�\Գ�x�'�׾}/���܆��B�վ�ϴ�y3�	��t��٪���^l��wW���۵k�ۭ�ۓ�/���+�W<̫�j߼ׄ�\�+,S��m�h0�$��a	t
����Վ�X� ˭C����2g��C�����V��� ���DIC~BY����u�	��?doz��Q�2m�g}���H
�Dو٘�0ԻjCx�w_����;r`+-��@��
2�0Q�͇������ݾ��x�f�r�����"��[��;���}p�}�����G��ѣ<���W������PiLt�a,����ѕٵ�Q� xq�>�w/(�	�ϲ�=\H�~E�p���z��7D�G�e%� ��G	%6n�/�@����q��f��쐍8'�*�̈́�H���@��|C�4~|R��%����p��fA����~S�/��k"�5͞���(����]Ŕ����ۜ�Q��n���5�}�}����Nc�b6�0����c0�H���\����7Ͻ�s���(<ok���[/��#+��ϴ/>��}����������)쇼\�O�_�|�}��v�ڝv�����7/,,��ť�!_<�՘u
ö0�R�ה/�\r3�C
H�_,�넛�P�DY@&���������7t-ÛD|�*��?��!�߅�T�.Ptƌh�¿ep��:���|K��=NAu䎤�{#��}����²�b�r	`��z�5y�j���ꚿ s�ֽv���v����Onn{ �,���J������3��YMR2x���)��ʡ�~'x�\�.w~���n�J�Xy�?�e��o���� ��˟����a�����N�����y2�}��d7���}`�L=�M��۫~;���Q���5G#q��32O`��cϺ�K����Q��(�l��|�B>���;��N���]�G)G�}������}�,����c���ϭ����~�ޖ���>8�>����v���vD�.��2�Y�2lo�|�~��?3|��㶺��M�������.�L�rK>a�5G� ��}2�׆��З�G�O��5h h�>�:9��1����0��feOs~6@��n���	��AnWaK�F��f!d72��X���(A�dԶ�R}Z�R5��L�"]��?�e����o�ܢ�����m��C�T��{�n��9�z�5nOP}�!=���>�Q��E���i++vmyzW\��B��=����j��
�:����>����o�&ю�����o���D��v��ڭp�\u9;���ɹ�:����0�?���z������9��M`�W#�n]n�輆��J����������&�K�j�mY�N&WϞ�1��N�Hڈ#��
O���~���O��[0^S92l[;y�`��S���]��D;q�@[������'�6ڍ���ߎ�l��mO���=�qeqYu�W)��b�l�%��`������n���\�V�x�S}#��;����;��x�u��SA5�0Q��o�q�~�v�&��� �dH9L��
	ZG��z����[�-��:�!q�@=v �^�g�ED��ԎQ�kR��������Ƨv�^�Lz�/��=�7n�o��l��L�����\;�3���{���K����z����b]��,�c��<3��E}��m���Z�L�rw�j��Xa�Q�4�B�����a��S�nu����'Aϧ��3�6�i��n��!3�dv�zEςJߍn:�hf�u�ՠ:ֻ����C�ߵ���/G�@�~{�.��޷���v.W��z�.�J����4�;·��d؉�ޛ!��*-+gT��ޒAʳ/ԾkmI����G�ŋgۧ�\h]:+��P[���}�=��Ӎv�������!�[7j�y�665��\Ȣ��E�Z�ߥ0�oU!��kǥ�o��zp��9^�m�o�@boĆ�f�OT��C#�3���B�Oiv5A4BbMl�//��wȟ�@6��1=�n�K֝ ��S�c���ݯ�JU�y��Ot�F�l�P�t�h(m�T�o�V
&:MGj��-���N��d�r_Ӿ}��֭~���t�����MM^|'����}������~�Y����ߵ���+M`�ۡ��ϦpK��3� �4�l�N�CL�w��*�7�WŃ�@��wǘTjB�IN��)Or~����U����Y��K�i�
�XP������6�1�z�l;!i��	d�t����v]w���B��*q��0j#<�Y��Q'��<���G�a:L��h�.a�W�5�P��$�ͫ_�5D}�t�/�IFMT��A��0��)�B
�i�,#�_��F%�ɤ����\|���ψ!ޤĎ�z�\�67�)z�>��>њ�?m�}��?���,CU9��k[���g���?�����w�ۣ������6?������󋲒%|�j��k��	��u���F�ftS�0��-�h�n/�b�HR�xLi0��u�h`7r��p�s��V�/�������s�����,~Ǥ2B�)x)H��=5��O��J��n��l�h�������+.x)3��>�/�'���N��e`llɡ��u��B�6?�Ù��j���)��n$B<�N�td:�8�FY��5�߱��z1D��u�6u]4�=�u��<L�IJ�B�	�=p,m&�X_�ѡg�HS���@z��ԩ��&����t����d���W�-,ηVd�*�> ��>�-X�D�d���n#��İ�ˋ�>���%��y#�pxpt�����_4�`�?�ЇK��V��S��W	��;�X�	�r�2M��5ce��t����I��·�n�T����m�z�J(B;:�HO�%zBҝ?��a7���$��}C>�����P0h�M�'z�����T�N5maȶ[>�Io����d�"&�C��X�ŝQi��W��"w\v��F9���8.' �����B~GU�zy��m@�J��E�\b|t�����<Ƹ���r);]g���<����"�pP����::�x׋[��Aެ���۱�K���3���}�է��_��|Q��ګv�����ڷ��j�}{�ݹ󸭯ÛW�r���ބ�����b��W�2 �
��Bk��:c���fS����;�4S<��=D�tN���a�W~%66����F><"vǒ��6�}��H�	�(N�4aE���B���ɯ���
^���Q�<�*�A��; G��bp{�e��4\Oh�l`����Y�O6��*���S�
���6w��o���*���3rH`��T،��6[�
;5�2�J�H��x䙻��2<a�;U���cO��䝬�45 y;٢�$W�����(�usHD�����Wu�W�gp&�����c�M$��w8���W=?����:���T�����a�+\$�C���c�R��rP 7y��$���A�YH����]\\
\���	�xqa�:��
(����񪭮�l/��2v1t1���w���bb��V�l[�#�\;: P\�C��>�h�V]����)ڃM�����[4�7y;�38ӘF����e��Ճ�Zudޡ�B��^��f�A����)����0�"�8���o+���nQ���!C\��Ba��Q�QoAI0&xL������p/�LE'���s'�jR�����,��^x�#\���c���c��>=�M�J����PG����N����+�h�C���#]�^�ԑ�@��3��r�9�� 4Y�u^
�t|�h���ި��"A0L���;]ƌO�YK=��L�����AB�w��V<eC��v�rTP�;g���o}D��O̭:�>�$��G��4�m>�jSٶ��6��c���O�˰����w_��>�Ў>�����7#��ݮ\}ھ���"�y��̳o��[��P��ڨ�mDy)PA�<���-��Yt!u��	����_�u����EZ��fDR�/m�UF�Y� �A�C�7T�Ƀ�Ҿ��j|E�~P2v�߁o�a���\���\��;ne��^�Ǹ-{-ڌX����O���ry��H5U4y���
&8�6y�~�m���4nO�<�Μ:e� S��R��MO�H��7�fb�I�^:�	�f��hEWf��>#?��?�+�Ip�"�,п$'Mt��evt^�Wy+��}Q��^����F�5�I�=���!Г�~�{�rH�F�κ����ڃ����[�﮶~�Dt�Q{�d-�������c퓏>h_}q�}��v��Q��WYۛ<9�N����,�/��1:7rRx�c��Z��_d�e�G���Ȯ4�	c�r ��L��H�uq�ޟh��.U�o�J���~f�b�����N��?a"��K�Y�i��۸ۂ=�6��{�ٗ���51̄��h��U��60��4��`�ꑀr+�Π���;���7%��^m����|S���|��&QN��c&Rz� �W�vh'����&�:���Xr���N�	�.=�&�L���e��>��� ���)��C�^?�U�U[^�kgN�1{�}����KϵS'������&����v���v��{�ʕ�ޱ%����[��>/�q�m<H�u�;ì[��'��-����@�uӅ�SQC������	�O��� �wh�,�]��P�AҸz�NI�"�Hsp��i�+(�|��7@g��]�|g�퀱X�G�&�n�܇�����x`���;���L3��3���{�=r&�_�\H��mrS��I>�k����+$׆���K~���g&qF!���a���/�@0ˈ��b�`׿�Q'���7�[.��M��dH�$��:��`�[�0�0�ï9�"a4bb���y�'T�n+��	j7�B"\Zfwѯs��썳K������o�[m}mCg�/���f�g^����wѷ�6�w[�C_�X�����2�@~u���4��u�/Z�O��Rݦ4?��fdR�ٗ8���\!U}P~��˘"��	��X�v��
'�`U�)���ޅ�4 �n|ޔ��-ɦ�=�\7��-���'�T{&�H��`�)xk�NAL�>8<2ƥ����Y�~(�n�UϦ��\��
9�������y0��*.�7b���@A�6Z����!��#i�qvDt@�;��t���
�&�e蒆Q;��Jk�v;y�@����~��O�GϷ�1l��6���ǯڍ��_�����^��f{��ցe��V�u�,��Bo� �\vr���?#G���@�t\*J0L�}�=@��v��b�,냬����B�+�T��K�.7Q���!� !�=�c��>�T����/��ն�e�u/�\y[�Ez�4��L����%����/AʼYu�,�- J�q[�n�����,�ʎ�m	�ǎ���B�� מ��- n�l"C�g�Ge��k���E��p0�)�=�21����-~�v@�`fY�w���ɢ� ���0�l�a��.K'��ŋM����;������{�޽���qӖչN�:�.^<�>��v���v��r[Zb��T�r��
�S�6�Q�U�XuN����a�^���3t\��Ua��_�]��ޔ�����DӔ������qw�(w��q��=��6C�	@L�Z�&���!��t\���.�3K��8� 〽��f���h�˫�i�ǉ�A䵶��R������=��Ν;)�������ʰ��N�<�,k���J�a����+W��c׮�n>i/״.Ȩ��{lmd	&�T��D^�۰�v6?�L(Uz~K�������!�Kػ����J�Eo����`d���u�	EΆ���s�e9#�g���,�S�7�`�V�XX�/��

I�\�aم����	�v��rg�3F��L��4����0!&�A�v@'�D���x�����4��k�~��}��θ�߸�=^�=T���)��R�A{��3���ζ�珴�Gٞ]S��?޴�(\֤��;�iܪD��n��TH����#��I�*�ׅN8c�tt!0+��`��Y�=�ա����+q���BQƬ�G��7��a?%X���ߧ~9�J0�
�zeܯUN��#0+z����G�P/W��ǳ�d�>lO��«��'ڧ�^��>��a;~�h[YZj��iZ��x�[ٮ]��~��ܛ���Gm}c��nk�������&E��\���r������)��8���9��80��o,��x������dѢ+��?p������JV����m�S%`��n�rz���E�0�����_ƭ=>���:0��2��ծ��p��&��R��ƨ0���/�[���@'�L�U�i|wp	.�x`ljR��������^���1w�=iW�ޖ���>|�ܓ��\�dw�}$��s�h�_vm��ۦ���I�,��j'��D�~���VR����?��t�}[xG�	�)y-�JtxT�E�d*ku�d�G�{�Г�FjQ������yW�E�z'�=�[gz7���u�jtU�[F�`q9y�mn��e�b�;����\��K���3���ޱ�:0\�d_x�`͸~�V{���%���٨���w�K��:�v ����a�Տ8�h��S�I��^@�$ÿepղ�3pg=D13Oa�O���0߁�`���	�C�!_��=�m	�P�}�6lӏ��)Ľ�t����3�,	a�w�=�3Δ�Q��z�l����y=Uyҋ��lmk����w�-,.�������!�/�����{��ﯷ�tΗ̞�\�E-paq�?��.^<پ����>jg��J��6֟�P�T9�T��.b�Y�Qm���
�&�Їw��&��Y"�j�{�\�=t<��K�����Yi���x�o�.��6z�����ʚ���'�[F� �{���)�n8�C5�._8]��9�9٧s%�	�3������f��9��6Ƴ2~�%�@h@��b����ꍶ��L�����="����S~���}Ԏ��}���������v�����7���7��;���]ޫ���,\r�~Й��s}y�A]�{P�dv3Ҟ�3L�$e��o���D��ϯK/�WXU�MD'@;��'�tg��?f*�] J�H{�m̂~"������|�<}eU���{�� ���,����<d��� 0���P�Q�w��F�0�ďW�r��p�C�M��2�|[(y���s����'T��C���'2��������R̲&�Ŷ)[��m�i^����;���g�������-��2�����'��k_~y�}����٣�����˶��\g�/U���%&�',��&߾��RXP�.�C�)CM0��U|#_�9�r&`ȿg�(w���:�,�'�A��C�G~��(�Ϫ+P�v 夷�!�㨫i}�$��a:?n�@�{�[�
��]��s�Ϳ�M�+�ǂ��O�����7��?�5^v�n�#�i�7��ژ�3ۉ��W���2���hf# �筃�Q�렲�y���v�g��V_v��u P����$x�(���ի�v��\;u�H�t�l���r5��>�./�y��ض��/�ݾ�LF-�j��mm���_��)��ȇ�B �=b)����^G]���ς>/�>�W��+tӂh����hծb%7}m�� a"�&�9��&�0��c ���m
�4P�L�@$�; df�_���gjm�����?@�]�øg��O�+u6!<��L��{i�7+���C�����6�r�'.u9��e�x�mL�(�2i��4*�L��@|�KeR���G6x�U��W��h��ĉ�^s� ep��d���Öz��t/��v
������4�GVcǫO�P���<�D�dNg�����gx�/�N�=�/�q�L}�b[Y^hK����W4��Ft����VW���ϟ�����Y �ʊ����7�F�aA��C脦�tl�$0;��'�]�#䓦��:@e���.�C�k�O�_�t%I��C�7�=�����DW�L���&��H0���AW�
�('pL�	1&g�D��O�asP�贠���5%s}�����U��%c���d�y�7�ϊ�v���M���̦78.' �<K@(y�Q���\FW���j���	��z���!n,(�S�c�PqI��,g@Ǐ?�vl$G��=e����L����0 *b�r]�����$�K.� �{�[l��Nٶ��q��Yݭ�U?@v�ԑ�ɧ��~�U���Oۇζc��%��޵��������=_ ����ڃ�O�˗�Jfa���c��Ƞy�����0�XF-k��F��!f��iEIz|L�.��ɋ^q�0r��De�.|����|�,6N�[�;[�IF�� �l��2^�-A�|�)�R�����.�ǡ�z���\���N����&e�0F��x��:�G.d�)�@g�S�R�L7@��#D�O��ۭ�jkCv�\;q�P;y�h;s�sq�v�P`AC}�B�H��@����4!B#�N��8�W�F��Q��3�5D:�!
����2x����g�S >c��Wa*���Z��'������]�qkB��2~�-���s�|��O۵�w�w�߈���yԞ>}�w�r�Ց�+탳�����>���?�=ƃd�5�;'r�H�A�;~v}hx�گ����ْ�p7��F���c��.�-!i�Z�2̏8Ӂ�=&�h똴�����:�XUt�i��$ޙ�u�T������r�{�X'�	���
�7��r{�	���L���ET�q�\�&��q�+O�6d��l��9��T�4����#�c)�b�؝1�����8Q�O����؊5�����si��	��~\������&������\;}�p���i���O�.�#��vN�4���ح[O�&hm��V�v����mmM���ɑ:�3���`Lv��6`�K��!��ڇA��s�q#8�=D5}�,�_R1GV��w�9���S����i`��e����~h8�F@ �8�i	C��#S���#��
��Ǌ7�YS΁&�������`k9��Af���sF�����`���9��B'�l���a5��K�Q���D�bb!��aP��W�(�~S�[�� �(G>�b��%>�k�j�"X��?<�@�n��h!��(O8ȝ`R�!�~ýRY�K띐�j�ׯr��
�C�y��C �[�mm���5/s:���Lv�
����on���5J��`�����c'�r�z�t�����{�f��Tx�i���08A���|o	��K5������;��!AX��� :��m�`1:���ա��?�H��*����Z���-���y��f��	�1���F� �eW;���@��1���
;�ߔA"���?"5��uf��i	^���G�
�1�d���txH�������簣�p���Ie�7�I��l�DY��̎��8]�O`��t���6��M8�]��a���-ϥ���������x�쳋�_��+����/]h�N�����Z�ń/�]���}�͝��?]i��p�ݾ�>_W��}�5��(��!lv�"�	�uH��.����◤U�!¡������Q��7���w�.�]-�V��)ޱŞ�>*�L
���[Qk�㶑��Զ�������]N�E��ƕ���'$�s2��~ ��ô�n;���ج��NG��n�y��������#�_(;y������h��jX�RS(}P��Z������G<���\�Sv�\�/�/~`?� O�l�B��I��&����<qf!�P���E�DS���$(�폨I��Y�8�B_�
�lC�I�!ǻ��A�4RF&��i��hy�-aK������p۪���r[Z\��|L���u���œ���IYj���i`�+���O����AVt;��#n��2�	��7l��2���-�|&�n�����ob��� Ɓ+a7��7m�� �}�#8�q�1Q.~\
tpL��]�>���Eq���ǛؼE1�/��o9߂�PW�^0p��!���ǛX�H�#��:]��U61��Ǣ!��y�ǑA����zSx0�������K��|w�+&��`��w��)���%��*��q��MX;��m�ַ�1�?�ܼ���v�d<C��W��|��ۓǏz���c���f�}�I��o	��ﾻ�n޺ߞ�)v��˖��!$T{��̺�a��Xc>�PAg��p,~A�OF�-��]^�ɢ�	��<�5W��N��I��t�a�'Qƻ_2��i~�$��ZG2n�c^j��ƭx�$�OG�;�Dt��2n��� �����XH�͸=q�q��[e(�vZ
�Ra�2((�^
pv#�! �(>�X*{0n5�H��#ϐ�.Du��/*�{�i����5����)� �2���ظ5�J*O�s*��l� ��!a��QZH���"�3D~�'E�iH�H��:�WE���/Z�;KR�'�Nm?�ݶa������&����/�,--�݈j�ƽX:�_\^�;/��u�k[�
��ҽGL�'�)ô�}X��tC�ޟ0Em�C7�Te��[F�?�O�iZ
���o7�:(��2dG]]�K]���/����[qQd毉ј��)6��D��T���L3�� �a ��e�1J��8tne*qڰ�q(vw�	��r�"�X��	]̂颦ɳ>]B�u���.� �s� �����L�f�� X`��l�֯���m`W�d�X�]}��.���M ���?!x���"�﷑P~�lyY�ِ���L�mccU��v;|d�]�p��淟�����}r��EVF����ܼ�}�ͭ����o�_�|�ݸq�=y�BK+�򂯨�
-���O��ʨ�5�4��ҡvjG׆�6aF�k�!*���MRdΫ�1�ff2,(1oWut�B �֭v	��i&r���1���ō�*���ٽ5��c^�a�Q:�V���a�W�U{d��l�sk��X&�����Hx�qK�&*6p�	n:���@jaH��c�����(#�J�
�;
Wv#�F�8"D���*KA���{�H�~*��3�=�;���k�.��t(e��;���_9�`ݪ�x�]��>^񵯭>��Y��v���o�������jǕ��v��������o�I��o>i�.�k'O�fS�V�P��4p���D�P�>N0#*�O)�$F�v��}1�O��������Ģ�cg�LL�G~
d���b̉#��9I�L+�����O�H'l̨�#]���D�H#��&��|,d#����� o����u���}ݵi��#N@�痄���3!q?� 0N���aQZW�d��`:�ʓ��_���<����q�mo��=����K��?��B�쳏4w_lΟmǏ�G0bx��铗����ڿ|s��x�N�s��ߠ��#��6v�̡�}���]a�|�9co����J���;��d��/�w���F��`�C4cRh
�=f�CdN���u'+fZ�I�5�,�钥���&���w��XԪT5���:�;~>u'>��1pp�߂�X�f2�r�K��qœ����:���8 ��08,���ޓLj��qfg�(�r8����?Q��ʴ�<%b:y�Rz�<�	'�B�1�0��;�Q�t �m	Tހ����'�����tf��6'�_���`p��d}m�������kmk{��8Ж�Ea����Y;��9�[����_�݀1\��<�.L��G��w�I�����M�o�jQv�4:	��A�����?�u��!��$�Fm���/�#�Ib��w4��'��d��`>r�͐o�5����ǁ�E�S`��,�l(sF	�4!�,��_���I��@'�,��(�w��2�E���M�Y�� �g$�-}��E�!��&�@kW)n�.����N�,fg��Rv�U.t���}f��hj��7E��!�O����z�`靸��hC�ܯ��oa���/�c���8qX����w���}������Y��� ���n%{�l�ݸ��}�����?��.�p�=x���6^ɦ]l�K+��E���֩W�~`�Ĭ�@����&������#C�y�qNE�75���H�0�%�a�'N�t��Q����V=��1D��~�	
�Nr�	���wPG����@Q����[%��e^e��~�Öc-#	��q�H>�Eyj;d��sk�ؔ�A�A.�"�x-���
A��/��(��~��e��.������P� �0��@H�5�͝
rbaHi�}�b�	I����O(<*b�&� �[1�#%��#Ë�o�ʅ�9�,�;�ذVC�`y����\tv�@�J��L �TG5���a��ӗ�E����0�6�Iv|�1Po�+(��cO���d]Ҧ��Gu2ν8:&&}��m��o	��0n_�5_�nCXX�}�<l��X�@���[��pٶ�8h�I]�����[шC���C��:���*N� O�4"�H�U.Ð�CG]b��qr��]A<�ό#jݥ�vt.ZXn@�G���n1�h���k�0������
A�3C��3�!J%�f�%�ǂ��l�0�Dh��C��*FZ�5�?I�8*�,�FL2L�c0�2	�r�r�"_H�|�^�D��t�;��[f�]A����[0�������$�H���~����Kuኘ�?�(��P��M!��-y�Xq������c����>>]ƥwle$xǶm�Ņ}���C��/>��}���6ryX���Zg��dخn�;���ﾻ�4� Ö�k[Z�4o��)�ּ�}��xu��E�^�z�&cP$`�Y} �ǡ=N2�g�Db���2����O��QV�9:�<�/�`Ưb�!R�`�(��;���Y��������0F�vRA�Fa#5�ֱ�֘�q�C2Ot�k�����s��2e^�<���7�;�;��OD;?�\&@�~agĺIܖ����+�6ly����'�ܥ��?����B�np�2a���ta�dA�nڸ�5�u�OѢ�u��{Ҷt��ŭ0�(b��FNeLT�r�c,�4lM�r��$�\�t��A`�u���[dr��萲�Lݙf�Ss"D�^�&W`�ǯkꕿ\�ʸB�(0ap�Q�(꩟���E����tHHq$_��aBɺ�"��u�[j_�w�ؖ���=�ʣA4���������_��\��=��e�H�W�r{Sd�2����1��)��\�.�lwf��a���������0!�-��T4N�C�zp��w�sE%�?�Ln�SU�Pm^��Vvᣱ�5`�eLs��l��;�N��7!Q�Ba1T�if0eu|��� &@ٿ@4cL�K�3' ��`&1Y�ff�
�Dw�E������*< ��t�|��}l�U�S0�m�i��0~�o�d�ei(Fh����gHR�u� ��̆�gw��+�'���蠬����?�	�U��s��������N��"B4�1q��7@�;k�����)7�-�V��&�f\�\���:ŭ��_}־���ѥ�2l��</��*>�<<vs�������?]i�/�n��?��m�����
�4��ƭ�K��
�{c�A2� J���:F��t.@eC��9��92�+�Œ?�dR����C��´�W'f��U'~ʃpdDJ�7�b*bMU[�qTl���M)�#ȕ(�� ?E�q+v���GAQ��y�z!���cI|��m%7�(��Er�����=d$�z22��5!:Y�H<��L"�h&vnѷN�0l�D{��o�����v��i4`*��13� ������'ªܘ6y�'�*�_H������Av�'H�Ԟ$I�1n�=��`��ޭ�b���A$�YY�0��2N#���S�e�"��'E��cNUZx�W�-�o}��_�0L�Sz����WthNr��ږ¼��O���o��>�������K��,�������}�>�dz��a�����%p���aX#Yv`p	��ݠ��cEBR�A�Y$��#~o�:���O#�v��ا	B<A8��K�����:�8A&��29�sԎ0Q~�\�"�9��g#�����y��L$)���rZV\�DX�0� ΂�,��A����N�_ͅ��>����п�{�.��N�A����As��"_2yW�@�b�w��������4�Y�T\����F��J*v�F�9}�]��wk?��l;q�H;x`�-���`ۻ�Vۏ?�m�w�]��Ύ-�]l*�+��[�^74?�G?���:��ܟ��|��&�$i�i���}���T(�' �>��arU���F��"��ܡOy%u�'��I�Q.c%2	��miD�}��V~�Ź<�:f>sSB��9o�0�]����\)�Q�9�GA$%M��f��f��d�b��vJ!��]��/�Qo!H�I�+����e�`_� E���E�2t��p*�c�D�n ��\�'��̴�@�4d�(/�|Y�_ǫXVT�@�DTtFwH��#F�7�hQG�[^鵍_F��ܲ܅���V��I��﮴?��J�r���5?���3���)��ϝig?8�:�0�6�|���3�<�T��vfRL�	��A^��~��>M�����I@���ۭ~�y��ߠ��!�d�X��%���0������α�x�zv�����h0���dx/O�,lI��0��0Q�ـv�'�J&�ćH���~ޙ����N��h�Co?��H� ����������=��t+��i2�I��Pq0�.-�<���gڅ�ڹN���%��d�֜Ϝ~�΋v��ޱ��۫��0l��)����5����)�G <�Y�n����	�i����.9 ���ը>-d'�vc�ݜ<���r�K�iF�u;`����t1�W0��k#a�ʏ�k,~�pwp��/�˲3�x
;:�t�V��ߴf�[N������a�	i/���7�Fh@1:2X���Wx̊��+��@%L�'��[9�&XH���nA�D���r��'��z#]j^�iA���������KS������;�����ѣ���.FR:�,����ׂϼ|_P�_g��B�~
�8�����H����&��n��A?�����C�v�*'ڱ�Ma5��f��H�n���4d�7�Pmdg�r��|+y�۰#�rN6���K�/7���L�τ���B�A�)�`FԻ���?{{���G��k�DzG�k�S�3!��y}`[s2����Xo~��W_(d'd�SY���+��Xi'N�l�N�lG�R��&�۰][�>^k׮��;l���j�~�V{��y��~L�qխ�L�T��FB�鯨	�vxK�'t�	�UhO3̿�0'N��E\r����@�zQH<X��Q��LiN龵�+�B��q�K�Q�?��7FR`��M��L�g@�)(�e:��	f�GD��j��o[��ہ^�u��<Q�It���������F~B&.��!�7���W-����@x�<v���0�9T�c�M�f��C�1 x��[����j��wXw0d����@���ڹ�)�'j��yؾ��j�F��O۽�����W��fk��M��|�����ʄhJ���ŏ���.`'k�'����dO��!u!݆�Ĥ5��ʶ����'��>��}���I�f�!�t��|ڵӗ��C����X�7 |@��L�ueGmU8f��C�g�g1t��Ah�Ř����ɫ��f<�!�'�G�Yt#i?b�qf��`2_F����wn�of�M�φ^E��M�Zu��?Yo�Q�&��M�ɶ���D�ZFŀ�;B�t�Z�mW0�^�鰎��?Ex".�j	�w�<t�:|�-p�S��fs�u{���ݹ�ھ�Q��7߷+W������
d��7'N����$�^e��qA	���Bag��M�%�w*�f�[�hG���p�w�/TI#����:k�։��Ĩ��Y�~��S�^C�Kl���L-DDd�u0��Q@���Q@�^�6`V� ��)���0K�]`���o��M5���;����f��CG���x��o�C����<�[�=!�������b��	G�b�������&�\a�J�&<vp�d��j��<o�o�i?\��~�Q���ǫڕ���w�������9� D{��i��|r���v�� �)��iص�	˓�`Ԃ�OC2�������V�⧏w����/H���z�/Y��Vz_��∜�0!�/	U~�D��1����?�N�Tq;���N���І]���.L�*�/�)^c�������\FǬ|V1����2W��ى��b9����b7���:g�I.\��Y���\����õv��#����o��7o�G���5^ᨼ|4ދN��X�Kt���R8�ς����gh�i����ɽ��
{툶�q���eH_�nM�����V��c���	~[�(�&�O��q03�п�D+�m�P!����j�lL�t���H�9��CbE�#�g��w�0`
M#oB��S��;F�Xq�P� g����=�2�i�S��@�j\�І���)<; �Kr��f�s�w���o�?�C��������w����"����?}�	��aޔ�ն�����@�	��P�]��a�8���2΀��z�������ʌ>��z��A띸0r��������
�Nn���`y���)H�	){�љ�ȭ����v2� 8�8=8l��z��k�d�p
������������M|폸�`���A�'9�C��r\���Fz�4_x�y|1�ԕv�°�\ڷ��4�,��1�-�8r���@�lD<z���?x�?�l�m�۷7d�>n����_~��EÌ��{�W����R��(ߐu˰�� �$P��gH��Y �����׻�B+b
��L��$�Q ;y�n�(�fab�z���w�r�^�S���i��X�R&s|�I@_����(�e,��)Gw0**�p�FЀ�l#ÎWcs���}�0�ʸ!e�ĨCo� i�d�NH��?ԙ�	��7�~��@K��S|Pv�3�
&��eκ���v���QL�
��E��&T��f3 ��1v>�ȸ�/_��y���e�/7��G�ڵ�w|i�����?^n���v������j���m
i����7�1�K��L�'N�$Ob��Io�a��?���a��}�����X��+���ƪ(��v4c�����8�=aV�-m�n������w���S�<�̩�Y~���$��l��$�;B_�8��A4�dŒ`A#o	�~��_0+n
��X��L�S�d`��,%���n�h���E؏��;��q����@���V�Ǒ���g ��7p��湵��v�΃v�ʭ�����7��j�����77��ؕ���Ç�������Ŷ���鞼◷#�|@�)AC�;�ә�:D�K��\W���$������C��c׮�ׁL���o�j�aP)�(�X�!bpCO�w/ǀZk|o@�Zw6�s�����R��. �<8I�g)�ĘL'�G��_�q3Mxz &��!�ʛ��g�6t6f�t��o���)�D���C��8�,��_��.,���q�^S$��Ii���I�z)�|W���`���H��@���=ߔ~�	/�� �x��g�A��E��\K�0h~~�����E5D�38�ϳ�����_8��I��#�cC�,�[ũ!�h�A9���2�l�&��P�A�ݿo^~G�=�|Θ�d�q�@X�ٽ+
����V_���i{���g���u�w�Wo��u�8H��s��M(7� 
�~j�nAOy_�4f"R�k7x�t�$x�ULD���9/ew�@h!t�rQ�a�����4�S����7%���0~G�rh�`T�@?�1j,�cSL�b����bO�n�0;+�QY����j��gy�u����
�/w"~��  )���q� �@�1�u��2D���8� ����~��w�^{A�@�5L��8��k�.M��F�u��6!���:w�؁uL�����Js|: �I}:r2'���䎮C:�*�5Xm��p`c}�=}�����nܸۮ^�ݮ]��n޸�=|�����檅��6��hu��H��o�L�Q�@�S�.(�쓪�ūN�X�ă�>+���
s�OOp~.��T�����"��r��0���*M}�u3���߂���b���:��Ӫ�<�(�e��(�L���0|���nڭM>��3C��������ͳ�� ����j䪬�q��O���>�	ِ^�	��#N���j{�m�>9ڔ�;��"�@��cn>^jQ_�+�N�8,/�]�gNkgN�h������^~*�t\��r]j�! ,�UtT�	F���a��5DY/t��d��2�����d>2n(#��yW��M8�
΀��):c"���x	��`Q�"{�
����K\�"if�`�L��&��x�v['>q���W�^�k�_��'OV��G2n���]����U�,�N��O��	s ;@daLR�_�@��<AFZ�}	�
���>�ӻ�J��P������{�ƈ����0v-��#DL/�^�7U���)d�@�[�;���2퐪g�#Q0+n 3�B��վc;��y�u�!>���:��0���v��E�s�΀0��]�L�ك/P�)p��Ҁ��2&ʮ�޿;0���v���^ܣߺ+9@��?��5��a,��:C��瘣"1 Y���FS�䇣"j�9Z�zsҼ�������v���I�z��۟�x�}�͕v��-�򋇃�_ah,ɰe�Vs��̖�yJ�ԃR�@�I����a��B�ز�q9.�Dx�#� bǸ!=��G7�ϐ6���T\�'�A�K�@_���1O�x�O�r��)����`�ٔ>�c�z�v`���7hCG�$�YP�GR�i��s� ^�� K��ڄ]D�������u3w�PVV���E�.B�qC���e�\ϯ [�3	U{�w�&�8,vC`2.�LB������3���<:,��G���*�o��a:�j�0���pxV��y*�_���d'vC~._��Z&���[��^�h�y���3O�Q���3�v�`G=��F#�n���+�Ŕ�09�o�i� �)@e��o��?���mJ��޾I$.��-PF����,�o����cpZϪܟ��@�穸�pRc
d}2�;?�n��U���ӈ#�Ǚ0P^�N ���L�= 󪌡-���~���N��E��Ԇ5(do�˘�̱U��L�.��%枍Zs�O��E��!
��G�'˯���������ڽ�ڝ��۽;�^���6�ݿ�9zQY攝��.3s2wv��u(f��G��BEk�$��Lङ� ��@�x*ΐ~K�6+$~�rз�9�X넰�8�Q�4�?X����!�'��1L�Y 
谏L_��yө��@�������R �����l˻�A�8��0Q�z�ۃ���y�wx��7DV)X�����5!mH�sG��;pM�.ci�f��qK�H��S(�
P��P!�wA`��M�g���@�A�YH�.X��~MB\V���^�Pe�g����D�U��Ď��0����_���,��?~��ې0��`&�6��*ݸ�����S�J��u��2g"��]p:�,����6�'��o�q��'b� #�=f��yЂ�v�d�o% �t�+t�3����p���f7�	(���1$�T{�����CқQ��u!�yW@-��Q�:�.L줽�-k�M�up�}ș��r����CRz�����4dz�cM�7<#��r��|�)w�mlH<�1p�|Т�]ǚCqG�����Hx(_f�*?)��es΋UdR_�<L<��q�`����3)�6B�
�ĚN���>�����,����HY��}@�M�9>tG��U	����鐡_�{�:9����Ʈ/�!��E�PZ}7�/¨ �v�eY?`R8�a�K�c������F��l�Ă_��Tgآ� ��2�@k��qq,���X�:�2�:@��Xi���1���^�7�� A_9��aw���;'r�yX(фK�����oU�Н_��\vm�a�� ��CYmg>9�q���Qxķ�g��u�=���A����ȵCw��,���̋rfa�O�P����9<�cVx��mݾ���?@�{_� ��կ�f���j�!�Co1�q��f��	,�p:��:�_�w�wtw��P�O������_`7��|K��PV�11�p���@>�@���'��4N���@/���C�ӝt�f�[S�;1Ң���W���(\X:�y��pE��Nc��_��\�͚Lf���ϱ����W:�8� Zxqk��M���~V�H7� r��"��p�T��h���a^X�ʆL��ZH�s�@�N ����r�����b���
H�F�9D8 ��k�rJ�r�J8YI(��Q�t�p@���m���*�[�[!Ȩ�5�N@�^�鰂����5����jWn�2�>st�&��q��%��Q��B0t��;�?�a�V�P`��ɘ)Pl������3iUG�Y�w\	M��)�=��N���	��ڨ����j���%w[z���/+����	�ez��^ƧΖk��� �'�w�!�� ��+?&!\ڐܴc�n[�A��Ա����ʛ���Е�Iԑ	]Z���p:=�	f��z?
K�v��*���z*O�)5#b���?�%��,,���]�	q�y
��=a��������*\Ї�K����{�:�m�0K>�0_�sx'`���i�V��B	0_��MFv)��l�О6�;�C�R�N��t�Txf�Y�4:��2#�縍�{j��[[��ܢ2�f�U�F?���X*�{����Q���;^慌���>=��Ǹ��=��<�n�$<�N����Xt��g&�r*'��z؁��M��0��t��R�`EJ@�g&�*�-~&�F��s�Qg�Ћ��K�2��>�q��I�F	�B�e2�s\��6��p�݅���<�d�_А6��˕����c�&�|PG���o;.����F��9�?DEm�p�%�h3�zZ.3�f5h�����6Ѝ���A�r�Ar3)E�A:k��i��'��64�m�v>������eyB�Ol�q�A��X��':��C��:����Z�'�h��Ɉ�[t��*& ���X[CQQ�Lѿ�z�q�L�;�V\�@�%GއE�ow��,�}�p��=��/��ĵ<�L���S�UQ.VP;�cQ�#l��I� @��E��`y����
Ii�`�2�������Á{*�����^c�:v8T�h����n<�t3��f�����M\f^���{��N켁%O��ڑ��g*o?�축ߘa��M��E�X��$�;�Y��G� �|ś�.�=���	�z�_4*�.a�-b�2ny��Mn[`Ƕ6+���7@�|�G��a��sp<������!=O6LO�Џ)�?��1.�N��%f��g��b����k�HSP����NrD8��W�RDg�
 2a�Q�q	䝄�-��*cblLA�e�4vfa:m�I�ʲ�ST��'9�A�~�ep��bܚ�0 �B��Jm��%f����@��;0A���_j��!Cк�v�%����<����%����;x��|���>EB������w|Lu>� ���0""z��8}>�e�B��7�E��'��{`�1�3Ť���OT��}�i���rs�'A���Lq�:�F"(�V?C�Qߙ6|}֜�s��q�,?�ƫV��O�&�K�f7@����d�.}e�w��9x���x��Q����+X�a;�	F]i,�o]f<,yo��]@�W��+�TG��Vd�g�dO]"�3(E�~?~FR���5�Y�^Q7�r\�}]���t�������?�l$L��`���~�r�����-�*U��#��zHV-�����};Ѽ+�0�����=RE�P��X*&���O�Q���2����"Z�+
oW�e�'�K���7�M>��ɷ\cZ v�u�_<�G|��_�HȊ�V����uƍ~FG�!uA�s������nQ6��c�6����ҝ���	#�r�"VY�A'�u#/���_4��j3�?2]�&Q�T<N�����?d���i1byF^�3툃^�*��%��C8�\n�v�m[��n����t��f������Y�><�
nH��1�		��YS�Ct� mn�FށF�+8o���T��������lq%U2��;F@�1V����?���T�hC�h�n�鰲���%���~W}�;����~��Ԏ���v
NE���udv�x�S�'_�M���3ow��B��B]�]��Ey���Q1����j��!�K��3$~�W�Vuu�$\Eޫ*��i⌹�Hg�2&��Q���U�D���Lw��/�t>�/�?�v:
=���t�g���I��G ?\��I���Wy�zM��	�ǐ�]}&O�E��4�m܆I'p�Bhh"O�x&����,�d6����n�]�n�	�>�����^2Ć��<�{� �\�3e�����0��3��s���"��9y�8H~v%��QN���E�᝔�C}�I�%�[tS��f��a����F�!'F>}�/���sB����R��~��}�%h�vC�	��D�!�wi��˒�<<\�
�Ҏ��#Z&3(�p���O�?��j�a3�k�_噄V��)�!�(����oǡ��J�0;�1�=�v8��F�d>��bt�?A�+�X��.��T�	O�;�^TDH˻H��o�A~Nh����o��5�}�Y�욛^u�B�D� ���B�SgQ7TF�;AD�U>�3���U�WPƓ�h=���6\	S��h�{D�N���r�B)�R���a~��P��w��}�y�Y�}C�LS��k*�ycz >�W����Ud��� yt�.>����!��=����̰���b�(9��';<��ˬ��U��^�,t�A��xu��\�*�u���0zM5vf�Act�B��8�C�_ ���K�5:���;��_���~Qo������ T�:&U�El��ř�)W���U����Agy�;���?�gO>1�ff�T~�D�\%��
l�Ui��<?��Q��:�M(y�?\���G~�*�����y� |��M'0�K�۱��ɓG�g��&0G�A�#�|���!��
 �\�HA�L�����1cJ��oE�dQ�ɣ�v��UF�H�<�5��f��(�L�����pzO($��h*m��,?��	NR���+��U���u:N����o�L螁>�1�X���>��#*�$U��L� h�A�Mm`�92h�?�v5^�N�3��� ��~	�l �r�P䇏w�;Z�G~���� 7;!��k�WB\x�O0Y�d/^��A/?�a��j@Ǳ8x�2*a�Y6yA�����W��sǌl�xR7�	^�}1��[�Y����З���i���D�}�?�SO�έ#�_��Ά����¡*[~��A%:�F��}s����'�m8�~;p�~�x��Z|�사��m	tQ�������� �>ھ�7�h�j��G��e�P&��Y�� ��̔�5�f!�N�<���N�$�.Ϭ)�X�F�6�c�l�h#�f�w�4��,�U�`\�/�$~YN��_�;�F����J�+�$��UY���'��3.�yR>��I��h�ߗ�03z̞c���\����>�%d��
.��X O��z�<$�������6�$!��sئ\�Sh����[�ېL2x�m�ݟ�on˸ߨ8�����]\�ި���|+π��W��q�?i�L��
G�]@�Bu�C�E���!h�_A��о�	�3ǐG�Y�H1� �c5A��!��\O���_��4��C���P�_�k,|�k�:�=�n�~��ǔ�NH��FS��0�Ȓ��w\0��IV���(?-�'�0�"w���m0U*FSȤ�I��e����9UG�7?g�yp��x�b��)a�]g	��v�a ��"���Ȅ��D�w�P��0�d�4,J��N��SeT�+
���wүC���;��{�@u���w��C/Y~��������(�\/h��\n���0�"�&I�� c!�:�U����V��l�r�/�g Ŏ��q3��"�����0yxq�p2��m&kM���#�^�n1�+�)mks�m��,ȿ�-..���-M�y�0����IF,J�3�Q�������W������B��y��y�iT~���������Q����+�����@��}U�C'�i��d��xL[��� w����f{8,��B��J�J
����)7�S���o��#}�F�8џ\V֯P��{�>J~�Q���LQrbTEZ,�xSJ�+�.�d0J`�2��1 #ɓaA�G�G?!�[b,O�G��tђ�����r�x�SH��_ry�8^F��e�
k��)e�����i�$��K�Hd����y��H�S}�,�|uSch�χ�1=��nQ�X�ܶ�.�<O��U=�}ޖ߻��=Ǟ���Y�S�S<lK�x�����[�Me�iG�����rC#�'���)��L����g���~t��
��b+�\r�y�͜��F�>.�p�qB=Ө��+�D%�21cN��s��ȉ#c,]#�?��c�e��N�td��n����d]�}F[�#R2�03��I�O\Hv?�G�W��k���3���1ȓv}����Fr�>5�:,�Ϯ��?���������w�S�&����G~W�t�EN �Ns��
c�!�����mey�;��Nm�99mܒL�G�
��	
�q��T��m����+{��A-})/~��.d���w�h�<ܚ�|��:%Ca<hABNB�O�q[��\1Rq�8�?X�.����vJѿ�_���&��V8�Wd�',��H��M�~��+0�I���0��q�6�1�t�[�B
>ĥ�5h�jK�ͯ��>&��u�J�	���'�n{{��5���~�<�9�@c$*�E�\��Y�D~��G��FA%��U�2`x�~/�;șƫ�e�r�9k7�|4I�{{�ŐI�1�1�m�)�Ә`�6D�$���s�W��'��(/;�2n�EA\b|Ra_6f�)�f�Ƙ�y�#ZL"O,��:�T�>�D��#!j
p�*���9��q4������!��0���T|.N@<A��E�zg�YP)�]\�Cm�n��|�xx@�_�-�Y�4 dH��Z��.A��	=�
,`�KY��W��rɍC��"�8QV�u�2��� ��3�xM�6�⬓�8��K���
;g䏈N���d���n��F���#9��o�9���"7�����N�6u`=(��+=�����za��7��Z��Zc�4�/��d�ul�1�CGx�(7�at7	��n�(�*<�N�N�l?$��#\�I�=���$��S��:h=00G�a�j0X5�u��4�����yiqq�-)l\^���Lxθ��Oy��V���91��vll��m=�����	��(��1Oh!�{��J�@�1C�~	'W��'�3��c$Ӵq�m��>J^ɯ[�I���2�1@_-�v�w�,>f\�{�q+:�C��R@�o�sY�`�x�����4n�-�d��o������y�,�xx�7컱j�i�b'gS�\��������s�G�l��*�}{,�:�����c1ggc�|�G�T=�5��
AE���)�XԷ%K���srP'���Xn�չa�e�c9�����M]A�Q�F���+#�	+kR�S@�O���5(��xW��?\'
u��1i�t�f�W�r`�,��P���C��2�L+��N-ןV\�~	�d9��b*`dʸ�G8�'����OΉ��UU:���x��d솠���5�kjB�GM��W��4ڜGLC_���W���N�zR��7:�+t�3G�Σ�ʵE�*9�D�?���T_bBQ"jN��˻�Z��!�����(��{�����PaB�ݤ��G��j��N�X��E��2+T�ҭK�����E#���� 0lk��d�%�y���u�U<1Ш�����)�I���KO\Ћ�DV�j+�a6ŗa�]*&n�jy-2��hO�(}�$����-�P1�)NZr�P�j��c-"��@H��'2Q>e3/��$ i�}6n�Gy�N�04��;b(]��ko$��E<ϟ�V��5'-���"��K}�u�з�ĩ�.�s'��ȡ��9�"��!1�) ����!(Ɣ_XO�#���,�ݢ�A�fŷ\������M7*e�x�j�@��eR�H��P�xG�6]I�5��?�>8�+qO7�+?�5;���#�/�;�[ʥ~����'^�!'F��P�ݱ?��)�\q5Q��K��m��I�B�Q:
�(�L'A���SP~�+t֌�H3�f�<��ϡ�r���!��X2f|��yh���*vU���> �Vj�|{A�=�u�3��YR6��R�\ tm��]�li��X����㪉M����@I�8���+��ju�,?�L6���e>#=���̑\!��>Nř#��|�Zm
��ƛT'	��![K���F��&yCB' ��k y-P�O�l�Qo�G[���}T5&;W ��C�aW8gS>�ȴ%��ʱ��^�τOZl���N2<��ݩ�+f�����6!�im��x.�^�|�?��>�t�}�ť����o�:(�+X��-������_�d�!�+�T�����u�m4^NN�-E�m�\z�h�(1e�:���Gƍ���j�\(j��J�P8L�%̰$�4��7���B�(�5�K�\��qk�DC�� ��c([XY+�����zPj��.�+�~�M����P}��IL�2�X��>,0�[2�^���\��$������|�H�,vb��8��şOoklX�<x3��B��������_\z�Ë��)���ɰEf�+������-�]76u��!��2ɺ��=��F�W[�+><�b�]y��p��bXQO��
A��v1
���.���.�t�q����:���c̱�+Y5��tR�:�zC�ԃ6��?ͅ�A� ���
���qK}10H��n�C��䪝cQ�F���ym�jB��"S/���H&�CtM�Q~�g���)c|�L��;��cc�u�2��YV׵`Z>�mIп���Jt;����>=�*y\�F,#����Aߡ e(��*�d�R�0������R�nKx0.7��#�X�H��	�f�(.��m&��j98�΢$�@�'�Xd��m����ƽK.2n{3�mb�ɸ啅�;�� �l����2�,�ǔM_����ɍ]}�����A;���c���z��a3N�S}�b������͘B�2l��9���B��2�= ;IO���+������V��K􍋮�+����Ejd$"�,���O��a�/�9r�y�;��.ɰb7vQ��/�]�_�ݽ�6����1N�G6D����d��|��ט�t�#;#wS��������!a�y�G�ǘ��Wd6��&�B�9�T�5՞H�ԏ~.㖂��N�/������e�����^�}���`��(^2n�Ӹݗ��GO��>��[wI*�����4׊��m�[+*�S ��ƭ'��8�6GG? %���m62�ݪ~�C�j)��q��@2X�'r-�ED�r�0��A�Φ��:XI 償��	�I��Z����u�
Ey1�2	ր��E`&G���J(�^ih3`�HA�ɂ�����2�sr%�/	?u��(&�>]Y�c4n�C�Tk��,��-�7�G�5��o+��Nv��G��Ǵ��8����8a���ԧ���᳾�VW�چ&��Z�0l�t���/�(gܶ8']aT/Ȑ]�K;nl��Ĩ��-
jcU�Q�����%�^e2�`�X�O��H���U�\MW*��;���e�C�������%s�˻�iK&&UB��g�T}X�Uo��M&v��dN��C���'�0�U�yM��Z��+.$���.*��	1A��е8
����b�~,��쪈����H�/�E_��y 9��&0�-�Sq�����'r!b��CԟQ��&Y��m/ԧ�x�W��� 8f6x�eGV~��_�a߾��@_c'��2.C�Ե��ns+������l�@���:�T1H�b�{;��3�s�O*cԫ�	sEA����޸��;��?����,�Azp�[����|Ck�l������v[>�1\�D9o��'ƣ����r�O�E
����J�p�5Ʀ��ȕǺ#W�6����+�?'�6nc�r��U_u��и|�2ne8�?W�\=b��C
k�<�̱��e���	�� ��&���@G��3=
\��Oe��*l7��{?�g��0����r����&7����+�Z���<�'�}[�|[YYlW��2����>阏�i �%sm�L���FU{��lblnl������1d7��&XW<�/iϟ���k2v�1�G�+�/�&�q�g�Ǭ��������x�x%��ƭ�|/���6[�ŃrS̚��c2n�)��b������yͤ�	9)��m~����ƭ��*ٕ���>����L�����H�yuN��3/��,�n1���}){7�vQ�;���M�%.K��(�Ώ�m,۸��z;B�(����$'.�r+!����=���Xyf�&a\�Ĥ�z6+�< �r⢣$Wqa_eG�K��G��qc I212��,��V>ʑ��`�w�h�j����3�L�!���uB&ur��M�����E�{d5=i�y!��&�����v�ġv���v��!��/��1�U>�s�e�ِ��� ޱ�##Ok����v�ޣ��ɋ���&8��d�������Y�)~Ֆ4�\Yh��ذ�OW��^�q�-�[�\C�r�k,����~Mr*T20��H0T�/,#�2b��D��ϓ�/����-d�\xAR�-܇���h^J��CGdB�O��J�p�kk[���g�ٳ��Kn�P�����Ů��O%�V;xh�<��X��#2�'��0�h+�7qga�B��!�t�(/�`�dmmC��A�pZ�e��U4U�I��p|�S�{�D�N�$�g}E�Pڸ�����
���A��;���.��1�|�g-�o� uآ���9�V���y�.8�R]�С�0p|R��A�����J�_�Q��Чs�y �\ys6��2��h��k�,�L䥏RޖN�0&��פ'�D?�:�߮~��ϯ��<)�dp>�I��K�j>�Zy��YiG����*�G&v�����l<����erpY�	o��8�R5ƇI��ؑ�ʂ�T�N��Ӹ�ξea����s���F-����W=ǉ��`�E�k 2@Ϳ��	G��Ć�d)�^;�vP�U(�y�(d�&`��G�И��TlX���\T���9����0f��u�A�Ɠ��j3�e�+,h>[��Ά��C�[h�..-��}��K;�ڸE�@=�ܲ��P�iKF��<�[۵�M�=a�nh�x�b�=a��6|u�����0eEaQO��ʚ��k4q�A�C>[���}�q�}�XX��S_`\3)���ֆ�-�n�.���q+]�r$ �q+�hkMƭO������y��!�E+?^�A��C^�<؁nz�#F|�1�ń�F�V��'m������?�_��P�2�X�r̓���A�Qh�tʸ]� U>W��\&��[)��Ru,����9�sT��b��8�����"��lp�CZي����j��-��\�@磑Ⲵ��o��Q��[�HB�D��� ���$PnuZ��U?�#/�S=ѱ�<�]�F�|a1/�Щ����V<u�n�,>Y��1����\J3�9��+9 �4�q�D-Z\�|�J�g�Z��O�
*=�p�L�E3�T���:�Q ��>+�9��;�j��eL��>:M<�dx�j�?8�.~x�}�����3���mE��;��3���Q�إE�?�D~)cxC}�ᣧ�ڵ�������{��UM��:M�L�����'�3����n�OoǏ����"��vߖ�Jex�䲻�kY�������j�v~Y�i{.����u�v�y�n�u�^[}�ܲ?v�}��v��i?A�������6�n}���ŁE�}S��G���+��͛wڃ{d�{ܗq�-C��S�[k��N�Ξh�ΝlG�Ĝ)n$֯�jK�3��t8O�[%���A&/��M����5��I{�P��d��[�BvH�h%/��;
��3���&`:<���3HE�a,++c
b�����e�����6?(����e���Li\!�ظڰ��8q*H	:�H`�`Tq²��ޞ>Q_{���+�iT�P1o"���s2�1�6�^H��s���Q'�p�vI�%��a�C�0mKZ�=�׵��x��mjp��}o��.2}F2�0�|��_>Q6|��<u�z�)��˻5�3��A�z�uE<ѳ�
��Q����b����:�dn��H\��ڒ���l�b�b �,/��lTxQ�9���|������8�z��gO��Š��\\"����7�$�[��0f��s҇��"���H[Қ��W���7k���I�T_�l��P���q"���+N�W��N~<oh� �҄@�/7���xG�]~�K(��!K��9]Bz��qkՁ9�\�v�����fZ���H�V8N8Y��0��C��\.:�"�9���:�>(�W�q�-#��M1C>�G�����$��[vc�����2nޔΟ˸}���N�_���f�Cl�gِ�|�)�-°� �;�l��C@7	zr�b�/vm�'1H����RR�[��r8��9�T�ʈ�q���5�-�(|Q6W�}"��?v�i$�ߴq��"�b��\>������(.�Ildb�v7����������Ӹ�p
a���	Ey�V��<ߒ�D(�J�ZXP$�����
°���ƭ:B�4nٽO�8sq���:�:��[d�[��or�nK0/)r�'Ide���k�V2ٸ!���b0@�"S��2<�q�$rA�1LY��,��s"#A�ͮ��E���⸠	2v@�τ��Gi�)\��IL�/kp�nX�������12b��K159r	�E����`��~u� t��@G�X��?3<�YoBYr�0��_�0���B$I'�essLHOۓG�4��o�~q�}��'�w��:��v�衶��U��6:Ԁ�*���Z���*q*�<<���w�ڝv�������i�c�c��}XȎ9�.^��}�х������?,n��#Kƭ��ҊT���&�!�<޽7eȍ�TC�&�۷��|s���ϗ۟��]{����g������g����cG�|�qǴZ]�q;��־v����O����w?��Wo�g����dXi�s�����2nXh��$��>l_~�a;u∤����ox՗�*���-�U�=s��I���d�=�A���]�Ӯ��:��X���KˇE��}��T]a��\�Q��T�L���:����.Eߌ��oB\�Ǹd쮯�����GVts�}���v���
��̃U@]�=��F.�"a��~(}�02/q��ɓ0�oߺ�v}֞�n(�.'�2��w��@�{Ű�h`�~eyы�!�a!.���a�!}%���
�/�I������#؜p������E�zb�,̿nK�|���wRG�M5�.������#����2�5`��K����&����rͧ��)Cc�ݹ��W|Ҫeܲ��J�����n{�9|��IG�?"�,K2N^1LtPA̭�)�J��'�w�<�����O_X�s:���_b�j���6nu�ͻW�$V���q CL�=W�:$#Wk���{�y��C�1W�s�e���I,��������3�h`H��E�s�X��7�n���P�w*���"�]~�]��i#���8�g����l�l���W����Iη�S�9���6v5rK,�vBc��Q�a��e�j�F/;�2p��¸�5D�=�0l�)㶐+�ܞ@������mK�/u�ɜD�����/u�I�ہѥ�<�
���C�#(e���|���Is� ��J��	į�[��c��r縲�H_mW��e�c�P_�Ԯ�pK�ʐ��0�[�@!Ȭx�n�;�e�*��[�s��$U^�q~9�2?䴎�w6#䧾�y�W2���x��@ٿ����2n�$�ʇ�@<�fZ�IY���@��~	�v�w��6n9k2`Jq���j8ӥ�����|������ظ�,�R� �����2n}k��DX�D9v��W������A��z��(�H3�3U�"�=�����|V�=D\z|f�zIO6,rv���X$�����bmM�L������ �X`���{F��1pY��{-�Ի$զ��<rFo�#��~�;S@�H;�Ǹ�/Jv���#�[�� 1э�۵���Z<�ڿ���������od�]��qpI}B�ƶX>]�CX�mh����&�;wWە�wdL^n�_�n���S0��m�z�����W���|�Y����N��e�-2���^l��R�6tu�,E����C�,:�p�]�H}-����7�?��w���/��E����>�����F2\j�N/�#����J~du�<>�٧���m��Wo<l�����x��~��&�g�{��{6��ֽSw������~����>o��>��a 8҂�%��r}�*�C�?�T4�=}�]���k�~w���O߆���lnbĬhB�E^��7�����q^I@,9��~eY�"@� ���֘d�i\m��=�'Om�~�a���~�.����)�⒢�Ԣ�2ҥ�l�fS�����(�1��������k:��}KF�S�6�-�����l��x��֥�&�v��:u��9s��;��\v����+Q����u/9�DxR�$Ύ8��<~��ݺu�ݸq�]�z�F�w蜓q�ue�;�_����'dD/�݊RK�FN���\Y��w��d8�_t�Y� u��9�°}��q��=�d^i��ܗ�!�Sk��gz�L?L*����v��ᅳj��:	�|K>v�i��o�.�Ü�r��f��+67���ۍ�w�Ç��}��T��!o�~�f��[�H��v8{�d;��?�t��>}һ��K+��V��	Cw��N?���OOdPݺ}�}���T[p��7�'1HM�vՄ�	���~�v�Z�k}��K�8���l��6�J��������r��8q�9	�B6y�-bǖ�8!8v��[��׉������c�s{H���%�(,���9�a���ot�^܊�q.ፍM�!/u��=�īV��A�e��WQ4qb�D���ˉ����Yܷ�`�R�4n��hd�p���d�э���[�p�s��[xз�d�P���3�i��vE.5���G`�򶄋��¸��R�|0��a��,f�a$���ƭ�WMR�%�9��J�q�@?�jL��b1 ��[+*��VvnV�ʁg�����[�(Y�W͒��
g��g���Y��[��[u.1������:�f.��cp@F��#G5�l+�q�eI�XDbW���E�vMF����:�.��Tg������. ��������侶A+�q�[�'(�:Bw�b�X.�������ux��/L��cB ���cN����kkO���74h������������q�T[d+��� �^
$�K�s)�/֗*�ݓ���֝�2lٽ��ņE�W&Fv�Μ>���?�}���n����m�./��4O��o����Z�h��G�A&�-n?Q?d���n���������m=jǎm_~�I�?���m��W�N-�_qR����\������.�~���������?����~h�=�r���!�X��}�����o��N&���v^a�M�w����ώU2i�إ�g�k�ƭ��nx��7۽�Oڳg��'-:��4ι� �(�m[��a*n�	Y�{�����>��"�{*i=J.�r��o����W��ڧ�o��7P*ƭ)�S��z�yu`�a��������u�����˷T�[�����|��x�׸�%#K�����k^زpZ�𢌩KϷ�>� ��t;q옌�%�E��c*��r�Q�d���Be�`!�}�A�z�V��������������.���H~�٥���/�����Vd�r2�W}\w��B��w��ǐQ���#���X_ cG�ZB�Sw�=�������N6o��x��/�Ru��g����W�����>���%��a�c�ǨpQ:���8x%CZm���������e��m��>�A�5�����8�R��S�B���7e�ͫ��O>��>��R�L�q�"�ed����)��?}-�[N6d�j0>�	�5���N4/_�<w�\�&,�$��[�xT�T5rV�ué����B�I;Fy8J�t��Z�q�H�I.�Vu�Z�6�������ϱk+[ �V'$���=r�����u�U_��e���%��܃WH�>��C��sX]��]zQ�~�u9]��������r静��.�mVi�a���и����:ɻw�Q�{��ǚ�h{6P� v�K�'z�"�1�B�@h���_,z�ַ%���=�[�5/�T�FC�1XF���B��%S��*ƭ\эj���
'�a܊N��vڸ����k�_��s_��@Y�@T4�#dV1���$eRORr=3E-�g��Xu|��:D6�)�r0��y� ����!~�+�"�w�p&�A6RUtݒ �p�|��L�M��r�ظ�U�T���A� ��~��5���j6^ ��dG�5`��çO�$|R�Йv��S�3'51�9#<y�4'O�e�S'��r��;vЗùL�}HLq?��t*����ǀ��<F��E)�1����|b�Q�����!��;ĉL���?�r���P��8B)O��1A^w�t�7׵�?���_liQ�t�d;&������m��-���t��ES�d�ck]��-,Z(H�p[�O���;><k/u��B��3�*|x���K�Ǐ�B��h�� v��Ag����*�#�qi�+��vۙ����Q�8Ѫ*�l[{�xC�s �۝;�l��Xi��G�1:|���;&�З=�q�PWt�!��x�<|�n�z��?�A�˱�p2(Qs��	�+�}�q���9-BG�Pقt�Q|%��B����VI� hܥT>"a;�?�xC �ˢ��Pq>v��h#O�t��R(�ߨ\ǈ5̳"��ת��uJ��2$ϟm_���=q�Z�ɪ$٨�W��Vlʡp~�]���ï�>![T�-ˀ=x��9d�=�|��6����$��?�ʏa��Ω�?�A��矴/et~���v�̱v�Т�̵	�����~pi����.�­ܟ~N���s��"�HF�^{�R�}Mm��sͅs���_^j}xZ��K����E_�8(#�����x
1>WT�d1J��!���iYq��� �=}�*��v{������d��f�{��̓'k����a��W��ϸ�\�t���v��bZ��d ��%P~NJ�����A�ɲ����m0�*Á1�ƕL\����[iHz�k�4>��\����l`s�����%��j-@��mE')K�3�js�<�y���0บ�[�dlI>��EƊ�46mؖAE_�KH�E/�^�?ͭ�9��B�%��y���у�s�̼�5'��s��N�� ��(�q՚��Y��r����ؑC�_܃{@m��9�����5>x[��4.(��r�t�8��Œt;��2Ŝƺ�3\=��yH�	f���� x^���}[5d�P|b��Nh*>�pt����UT]��	 �����΍����V0�i�Fr���*��������z�k^�P�	��x�E�g�����r\^�c~7��[V����|�k�N���蘃��� '��k�c�?vȶ}f�����`ܚ�)����J�(/&�m�J�V�\gS��T/4���'y���s&�[��\4sq��[%�2i2�]xW���Ɇm�2l1j9S}��ūL����T� �pY��}p��ǰ={��=���Nb��i���hg�>�����%�|)�o���C�;�=w�XY�d�q+I�,L�hԎq	Eqeq�S܈(,(��x��>
�n>�i"!�c\�*��6�w��j,�naܮ>���.�c����s'��x�����:��P{��i��κ����zw��C���"|�V}	\�A?�'���.jfV����d���X��]����S��k�ς�������!0��?y��=zD��*�Y�w/�x��W�k!$@�Ka�ã�����֭'�ڵ�r�� }�˳\���3��Cv�ym'^�R�%��1�S���������6l��������~9I��=&M�q-���L]�pF�&~�o�X����+�<����&x0�3߯��x��]�q%�{��]$�-���K\��K�����l�j7�A&=O� �o�"\<B����\C�1l6d�,j�R[�dFxJ�[��9���������L�(����P��%�t1L�>�k��)-��H母�gO�I���s]y��/�U�K��파��>:�>S�p��hP�@ҸǠf�Ɔ��4�x0���4��F���Y��kjǗ/^H�m�-�6@�����ܱ��6j��2%� �ڍz���,TRȧ4-	v�ƌ?����뱣z��M�ׇ�C�ݿY��=���/d؃���x;�yqY��z?s\�Y�����1����U�Z��?���|���d��/`��ϿҜ+�o�||����Gxs��d�}PW��%�$a�j߳-�l�y�8�쬕�T��ωs7���֜�>r �:&���0}�_�Cd�(uH��`��m	!I�۬)���������o��aˆ�"�ոbז[����:�=�\��>�[a����<=��#���?���C�[��M�Z2q�'�&�K������Yk=���G�8��2,c�Um#�Dk�Q(f��F��[�!����#���t�� t�d�Mc#Rh���sW~c��F�|ծC(~q�<x!�(W"q0��1�eP��m�%�%w�Ϩc�0&�;�[lE����\o[j�y��˸='㶶�)�FlV�7nc4�R�0{���j�i>6Hm��T��wn'+��$C��ae�\J�X�
��%�U�Q���@ee~��!d�V y-�q����O��vl�����eMX�t��N���6����A�������ǎh0˨�P��"�P�YAՍ����L�[� y��w��i`B��C��u�S.�K�ܢ#���c��_ct�X�HO/0t~��J>c���<!�B
��ԁ�EE	
V{��D�r����>D��OK�'T�-��6m�~��7��!��|�}��o��p�����k����_m�/s��h��ߘ�e/t�"(C��P
g��/��z�Ev�F奋��9��#:!Ar��Ř�|?��õ�ͷ?Jʼ�~��v�z��n�$�����\kW��*�ڝvEx���v�*Z=���Ds���Ív��}�����L܆�֞>y$C����'�#&o��%�Ű}��L�|^*G���2�߶q�\F)�9:`̸o�'j<�w^�>sJ�L?��K�O�r���v��}����BN*�Ȁ>�U��?������������6��u���������W�;�:s&�#�!d�k�E<cb��s�k:9����v\�X�̚�'y�~�'�#�����(ܣ�RF/�k��!@��Q�)��Ʈc���7E����7(�I�y��m�b�}����?�fY����k��2�:�M�[/�9ˍj3�0emxj*�>�e�Q����5�(>y*��F�/>����aɮ$/ه<e����c�{�B�ܭ@���1�]zZ}��[T�^�����z���
q�Ա����������o?���<�� � ��w��GUov�1���}����1�V�;F;|��a��'�y�(��<L&-ʰ]h.��N���ݗ������y!s�!K9�9��������#S��O��x[ �բN�5y���mj�&���Z�c,P���r�H��,�\��/��&v����! �G�HE�4� p��U̼�l~����|^i���>*c������)��'�j�Ѽr���6<Y�ة�d	=Q&�+o��.���1�<�#M�i��o������J<���4_5���[#l8���'Ur3����թ��;m��}��N�N�u~񩾑q��F$�h��eP�(�Lm)]ۦ�2n��p&��0.>&��!��b�B2a�R6��gD�0���'������Y�0n��"��6d�����B7Hfx#@T,�#.�q!��R(��v!�e	��GʞڹE0��o���!�BF�(^6n}y�z�l�2��Q�l�k��-��H*ٌc8�#
���q��,����:I�a{X�:g�|nA`A� :�A�%�#���eQ(��xC���p81�b��2���{�V40�ts�3O�ܒ�a㯻`(�{ ?QT��):0���QzK����*�8B�<��hƾ0��{[���gOU��,|��F���`���w۟�rY���Ï�ۍ[���G��w���;w�}�O�>����.3����'K޹�ܓ���c�עʿ(���Aw{".���ᯫ��ˠ�.���Ի6*�I.\a���o/xhy�%�;�V�>3]����+-�|h�>�D�\k/^ʸ}*�j!\�I���V�p���ź�M�?sM�ݖN��w���`��������W����e����N�������Q�[���+W�o�����M�������w�J߷����j��@,���(��:3�:�g�{����_{�%Zzv��l V�c5�q���dJ\�0�˭�ài߃�.}.x<�\���1F�em��|�'�͕�{��?b���w�q<|�y.�?W�����z��W�ܒ�J1�5^����m��T�k�d|��~k�2�x����ڙ���9�>^o�p����{:�K�R_�����lU2�K����S��w�Pv,���>hk�w���Nʿ���v^z�r:r�i~��+w��w{וM���@es��n�? >��=z�b�{�W�?���.ޤ�o��j*l�t"��辐����|�f ���V�B��s��
�L>y�=y�^�}�A�3��z���̱��K�L�ܞ�������R���v��1��~ŭ�}��c���Ö+H����uB��l��p�Da��ٔ�X�! �{��sb,�[E��k�����®�tz��v��&��[2D/,�<O���\ҁ�SC� ��k�
��-�3q{�>W�5��:�|����4g��I�I�#�u�t\q�ڱÇ}Ց���=g-�ZƤ˒���F�Y�B
�%C�O^ꇉ�f�8c�޷.h���(O�=�⠵��dL:��Nٕ���}Û��Jc$�,�<q;��h��mm $���|C�4�a�2n���RU�}7
s�r�	c>B?�/�G��
����j�t�2�$�H/q�9}"d�I��~�su�{S:ꁎ��hN\��-W�Ϩ�;S;�4�����D|
˱�8!�`<�	�z�aK�@�-4��c��*WG�
:רrʟ򄁋��#�|�Y2F���B���d^�t�����;��Y�.D'V
uaj����g���}Oա��v���vA����%�/�5�`=�[|��I3��QN��1����Y���\�a`�`D�ujr>,����{�3P�P��]\���K���3�P
5%C��Qg8Ꮓ=rk��W@�$:�&��e S�����O�A�|��9���.޻ʓ����{<����.ˈ�!#��U-ϴ�q� O�?y�E���'Od�i2�l���W<��@}U�!�fy�������).���:q9{�W5?yͽ�W�=h��z�*C���u?�����;y,�,�~��_�����G,ʼ�i3q]�ݚ��	ֵR�/����F�Nq���3+2p5�������.>jd��u��q���?_n�}K��s/�6�k��Έ��?�%�UK��#K���32*N�>9.�2��p��[��������72�l�d�������]�ή\�%�ȿ%c�aVZ�e1��7� '}�̵�~���0l6�s���k��O�˕�5w �1���I.}G\��=�ws�O I�h{%H���/t�0�Ns	�I�C�r����-�(�ӟ~h�ˏ��o��W�H�|��]���]����vU��q�rq�sIcԣE��"ʃ}��ݿ��=_]�nN�<�~��O�o�������.Wu�eD��˗������J�㟮�o/�m�o��o�ﾻ���;:�zd�onqYF�����o'`~��m^�z�)y��$�i������K�^���E�F��-��;�����S���N':�urw�]����V�R�w��4Z��o���^��~�@c���y[�����S��qr���9:~�`�P}Ò{]O�I�t@{�i��:����x@����n�����>�<��k\Y�g�������Zc�gI����p��'��߭�'8�8�I���_�;���W�F��*O'��s\!����,�������<������pv	1���W�	uI�8��\��5���6Nd8ы5�����N`��L+�:��j er��O�Ht|d�� d[F��y�Lg���nh��[\N��ڨ���K���Μ�
f���ؔ���ڦ�j,�����]f��'�c;�q?r���'4e@�G��+�m�zNx��|ٻ��O���:�)����K�w�#�*�_�;�F+��*m�cH��x���ɯ�Y+<��d��(r���W�>�yľ*҃���sk�O�6�x�I���sK_���ې�̶Eă2�Ӫ}ȿ�u��P٤�C��};�Ɲ��0,84ZN�Y*���ј�
�7��B���L���;��+�y��2�VT5#��H�'����'~�(e�GF�uǰ�%|��d�k����@Fs0�2>�T���������~�s����v��_j���L޷ h!<vTƀ�J����h��o������(��"$�JF��lS��2p�������,�5F5�W��9��5g�Kp����\���R\��I�> �tP�e_k�Ykk�:���s��[v�H�'
�N�5yI^7"RU֬�U�5���Zݏ5U�9U��Jj�t']kA����a�}�'yoDtd���6��`Pll��D�|��)U�Pn�V75pH�|>�������1VG(����h��R�J���
��9r'>�af�6w��[�7��}J�ٴ�:�K�QnϨ�S�Q����Q&��3��X�y� ���i>��٦�"�l������}��0�5*�|��s�|�ǖ	�*k�~���z�l��U)�kYu��;�(�>�|�/)�lx�d��p��R�Tk���ͨ�S�r��\����)��N�n��(���O	_IIy��{�,J��k��R��R��V�R����c����<�}�-%t�L�P0����e�/��j�Ԅz$X�1ڮے�Յ�7ګ�a?�X�����8,��f�j�B'm��nn,K�>���P�	'�>�Ҽ���/g���>,?<|�/�Y�f5wF�a��T�����O�X��W�c�"�Ăvj��K�D���V.����_�*�n^v_�ǥ��Da^�(�f��a�e|��K)�o�+�o����*��y3/�.Y�(����Ul�`E�[[�����2�vƃީ��g��R;%^-tO�^�z+E�y���~P}x�v0k���#�nR��@&<������������ہ8�i�i�8u�\�b��5��(zF���p|�[o��gY��Ȋ�������*/���M�UyOh*�������	ŇR9�����j�+���+R�>�����X#?�=䉢��L
�P�.Ϥ���Zt�&-���F���9_�󊛕⺍�~���L:��da��o9��V�#�������h�TPY�x&i�!�9���b�i����x(���q<���m�gH}�!��c�ҹ���Ÿx|��M.����!�I���h���kZ�;�����1v@3�lˤ�K��QQ��
5r!�d�ǰc��=~�L��n����sC���[�`̤�P��!U3nHC@i��@��f>�k=�gM?��WIQQ&�}��(���FfQ� <���vV[�`����h�_�����LR?f)�5��M}����zr�oj;�[�v}���8������0��J��;��1��:W��𣄪��ņh��	�B��!�rh�r^$�T6��`4�d?����(�7����-��$v��Pj�e�"��p��ƙ2������Gy6�+K^��x[���à`�|zp�TZLpcֆ���OQzбhV�2�c�
�8�՝�����t�҅���t�8��8^�2��(�!�n�`�{v���]� t3�:�(�jcKH��8 ���zmLC�����2z�X?���p���:c��6z�J/
������O����G-Q�4�Q�~�'
Y���- 8b?)z_�	����j�A>��xV@�h6��m!G��+|X�1Fh:���3�f��׊|�1Hx��6|�V�gV�_��? ����JN*�#��%3$*�W; g�8̽��A�p��;��ʢ�X�_��)C����h?Z�vH�yS~��a���������So�祜k@T����vF�^Pڝ6He��U��3��X��"%��D����@=���uQ��^�k0PZή&�¹b��e(?�(v�X�+˚T�:�m%(t(�(q�_ۢ܄/^�H�zU~/%�_�m�^�x�bJJ�Z����d�W����ׄp��|�-� ET��Î��۹�������K�tRiI��B��["Zd�
ߓ��>��>~!�UMH4�b|#�l�P|1E\���.ܑ�}�dJ��mqiIt����gjOO�r��K��JJ�)����L���g���2�fZ|N+�s����<ۆP�<�:�V��P�[�ƕ�#�w���������1����巿�AJ����J�O}��?<)�}��|������/����?�ǿ����r���f4	cKu�{�Uo����_L�8n	e��l��[	\<�hB�^�?�.���I���|_�E���?(�|�X�>.�}�D����ģx����^a~[���;��$�+P��{>v��u���NS�>����K�v3��. "$R�L��@�Q�w6e�52�}�DpT��#��铚�iL̓��Vn�c��֓LQ�� �Wk��eR��=н� ���/�v`�r��Sh�t�(W�kq>?��}����w���:BZġ�]N� E��X��GQI4����!�X�S-�g�~~�`�8��pH����0 �5N���/���J��)�S�ÎS`�c_�s�-�	����XD!b������������`*����`�U�V��42}Yi�x��Nď��̘�Q!��x@��4������s��1o=�xNJ�����&O��#�Þ�2��Z�W��t*Dz-�j#m�>��i�R��n�a��W���ɭV��X��q ��:p�UQh�]��k�S"�h@��g��� �ƫ��ڃ�ʣ�&"�E��Qy��mM���D��r*�]n���u��}{;3[&5Ⱦ�ɇO\���V6��j U
�9�)���I_��Ӟ�Ȋk�~1ҹ�g�7�g�Lx��Y�я0u�����:�BU��D�U|)"���N���t&�e���J)���dj�
MS����Q�(�j
��,��@I����a) ���  ��IDAT#*��1�Ci�ć�I.,�*3og˲�
>�$I���"��g���`x��ã�eC
���x�+(e�crm�o�b/�a>T`����CЦ$�PŁ�7���hBi$Oq���0)^l�`eE��փR���&w.XY�F�����҄���¹�d�)  ���Cr�'y���lX���������q�q��y�������WY9?�[��·�������2�v���]+o�=�[�X/��H�/���J7b�)ɕ��5)��eymA����Բ�{S����X9q�A��S����g�d���#RV9ct�,-r�ȴx�\i�Z#��z�v��s5/G�'x��-H���sRnɏ�'S�H��^g�����z7?�~�y)ٜ)�XyX�=��	oY�P��2y�9��p�2{`Y�B���٭�}*O���NYX���b��{�|�[/^�����$����yV��s�>��^+���o��B��&<���O����ޱP����^D��P!������3a������1���BM�ҩm���1�6�q���?��>o�Nj�<�o��Z�-���9I���	�>ן
���/��H8ۘ\3~3�d�C^�(�ĉ	/ ��g���b�K���r�P�{/���$��{����
���~��ށ���F�	KZ5]�p��Q�bu��n�V��S*�I1	zpM{wq�'�m^"����m�U�Ǆ���J�D��<"8�����2ld9���c��HO�wR���2��l����k<+e�s�����9��aO�a5�z��S����H��V���A�@ab d/#���=1q����}��._�+u�	)�\���� f�(��D]n���ǿ��E�7,���Z�;�{��'ʱ��y�B+ޤ��z�jFU7�|�Ñ��+4�Иܤt�c���S�c��ʉˍ-V��ޔ���Di"����|E�+�	#��b��w�/���� �PJW���g=�PƔ��eH��>'�>85�h?���I���2R�r[FiEy���Э2f��<�'(k-B>&5�!��#�r�/��Ry���0��E��[�VV�H�:��3Ѥ��u�8��-^�����<��:W2�a[	׳�lށ��r�Ǧ��t��]J��Rِ"�"t��[��5�hn�T8���
nhuіYe��O�<�eum���hw���@�?�~��ָ��_�p��r�b�MH(�үū��(s_��jnT�����s��ؤ�r���9�=j�L�6U׹啕t�[��~o��8W�?��=�,�RT�:��[u��s�&�\����=�P��>6�-�mUuy�?5R�\;Y������E���?U��?�M����o������?�_U��o^>����Ө)J���i)�s.V��3�G��<�}���K�������By�d�<x<+�*O����|��_����	�bOE�:xH���CcV���۷�`;��̵�\p!Tm��1�f�t�~bT�����}R�7%7�?-+��*�����)�Se�5G�A"�sv�&{#I�Wh9�屔����ܿ�}y)%��|�\�9�<9��,&��rߍYΪ����@���zS1�Ǐ�4��U�ob���>ǎ1��D�&6'��;�(�l�Q����m���S�wlbu�����%gϰ@tRy��kN�88q\D`�`)� @�O-��ՅZ�4�S����Dp��ךW����e��A�*����i��~B|��'��X8J嶍D�N�����	̿~2#�_�܇�U��k�lxe ��y��U6���tVF�usE*�ì�r�:{?��������a�i���w�of����·C�����>0�i� bGN�uJ����Ҍ���3R��z�g�r�.#pf%g_r�K]�u�-Q��-1�{���A#�Ʋ_�a�6��ir���Q����d򕽩���ĥ�Ġ�GVR��9��c����(�(��	V ����)W�W�� PO��1wd�>�mJ#B�XyDA�
Q�]�X�C��N1������fm�7�A@��d|[t����g��@}	Y�7B"�p���{v��F���5,�.7=����Qp2��҆�ΫJ��m���	��V+���.K9Ji��\�=���g)_��l	77��1E�=�*�X�Y�J����dۆ[�?��з��A�o�r�^{Pʽ&U����l���U���
/ǝ�#�H��$���=�L�TG7��E�̈������N��;.�PpZ۱W`y��~aC��]@�}[<xQ���I�������Ϥ�My�4����eo4�)>n�2��2܏?~d��>{LJ�r����ŗ7���I�ꗷ˯uW�i��̯��՝�嗟�;w���7.�s�8T�����a>&A�'��M��#L�W<�V
��r�{�*�./�NG��S��kG<�����avS�}M���ت^P�T�e�=a�tj�?6�������Oޖ�6��xU���E�w�쩩����bK������$Q�αe��Z����̈́�훲8?_���Pu�W�*)�Q��q�7eNe_����J��6�u�m01U����{��/�)��DŖ��ƅ2�xÛL�B}F� 2���བྷ� 6,e�mں۷�e�������x��hM�XH��-c�dР�2�m��p�q����h�-��sc�s�˙�"��䳧����'��=���c嶉䈽D����9c�f�k��q�F�l���e��m�~ ���J�����,^a��U�M���TO���[�59&OD��dJKQ,�2P�5]A�ǟjق��6Vq*2֕���#�r��(+΋;�s�Cƾ.u� �>���FY��#��{`�k�F���$6�> ޏ�P~;�m곕�LA(pj�P�BF�Rb���g�9+
<����"�H֮%�-�z��Dxב&i3�s�P9�:B=9���С!�����2ql���0��uK��6�ɑ��ӿ-�Ù�{�:�tk;���`��  �jQ�hLP��%.H���p���T��Rɢ��51ϑ�h��aV7}Ӑ�tt�����z�o#��ol��r��.)��R\���E)esm�l���ޱon.��X�E)�r+�;��������	#��J6������B*�[B�����	Ӗ����U�?��I� �O�'âB1��PV��moz�eZL�` � uy����Z#Y[�����8_����-NYX����~��o�)���o|���WӚ�mI���LJ���
M�?IJi!!&�G'��З_�-�,����u�w���˯>-_|z����r�y�B�v�|�z���s������'W��⏴n~rMJ�)o��.n�sE�cQ��.�s���)��?._�@J����1�;�
g
�؎��'��L>����2��l�Z���?(eL�ɢaZV��]��,�΁�#��]^���"�����|:Ŀ��w��{P�{Q�&�ˊ۝><$9.c�����)OlաQ?5��e�O
�˗?�Q$*���,\NM���K`S�f:!���uR&n��_@��cQ���U�W�����1�pN�D]�=y�c��&��'�DG{��y���|���9k�I�D��G1���7.�`�+ӧ����'���֘P�<B����VrM>�ПM'��ɟ	�/����~H�f��K=p��GyƸF �Z��~PG*��*A�	��H�N=P��8�#u��Ӹ�������ɏ�.2R����3�=��'.bҘ�A�(�2a�}��_oH!�-������ֱS����ɘ�1�cc�"���(��_��3`��~����ܕF]-�V�!�.��r��T��+�Qv9��o� �����a��e"���sb�W�]�!P�ֺ��4k�l��s��<�Qe̖�"�9*�(�u�̡�+�L�Ӂ�qW.��9�}�M�K��X*�ȗ�O�8�C�9����3>i�굳��rV���r�&C�P���x2��Y�眆����֓�6ð���HBV�m�I�+�ado����w�vd�L���!�pVj��Q<~�|����6��O� sD�Y�u�$_�rSM��SG<'��BnR��S�T� 5� O����C*�Cr?̓�4����0��&���LU�O,�:��ǚ��C�QO%y��:D�>'� �B�����&j�=�g�!x���0����U2���? ͎�8�=�W�e'�_���\�$���(�*+�q3`Ч���ڕ���~�E��;�U.7�5�_\s<Q���܇{����ɭK���n�Ϥ�޼u�G�qf3�sw>��j�͍����ty,�|�l�pg����B�y��9��\�l��mKʸ&�gO���N����Ç����y�-�����:osԟ�>s-n��_q!�d��yyp�ey��My3�X�Q�Q�r�h��Tg&z\߻!�ճ1�#�˥K5��/'N�(\"�������g*3���4eP�Z�0�:&��)�՚��}tr�ɰ���}��↸EoS81���ܾ9�-q���ʧ'l&PiW�|�C7?*����-�؝`<{ےx�{��#����ϸx��L���LPpUT��*烈y�@�'��	Tg����N�f (��R7dȭϣ7@��	N2��:�����'qd�QB.�/�_�Gr%�(���d�?#N �Ddj��1�M�x@�ǌ�O�3N����4���%+�u�iu]Ლ�BC�����E'�\����VQqVTD�Ňd4\�ݧ���#�N�YG��c-n;��c8,p��@R���=��K�Yu�uP��+L�_Ǐ�����
%DY�%���=����Rp�z{�#��˟�D��B��6!�DA�W<w���k�aN�7�'�i�1V��tZʣ�;��2_M���,CqcUkc���z>���$��:���x���:��[7��3)�0;��Qu���#'���'����?�*�������W�����;嫯n�_��v��/��n�\���7����L���^��Ly��G�%�W?��c�i �P�S�!��k��ߺS�1�+����!heL���"��M�d��B���ד BVq�ڄ�2d��j�VҰr�+�U��e	/��#]\*뫫^1E��q�R��ӛ��n�/?�U~��'�/o�_��n��/>-��|��;�r����Ϥ0}q�z���U�w�k��O���������'�����=	9{��0Lp�H��uV��EYX$���p5�I��c�87�����.w�I�4�(�G�*�Y��6&d�GQ$D�[���/{a��)/&Pl��X��V#g�.�,�ZfVr��~L����'ys}�d�V�5V���2��F����*X�NO�=�"7�vs���r�����gw%��������!���K�i1.c�r���Q.	9U>�{Mm����Vn�D�=�r�"?��=� 7�z��z1�#��ښ\6ś�3���nl��/XU<&�LfW��h)����2}�|����۷��3g���Òm�������s��BY�L�7��f������Qf�C
�̛�����z�lnS�iRl�HC1H��hu�}�3e}mA�-�z�|����o���ꗿ��ۊ u��p�J�%:�!���)LԀ�Z���D��:H�o��ى��L�>"��������z$�@鯄(ul��oR������ǎ��QZ��1Gu:�@��������1 �t;W���W1�R���3�o�>�8��c�0�	1��ݪ��O}!	��ѿr���IV�w���'�~��"M�c@�l(7�`:a�2U����BX�m�&�[�*��]O�~�SQ�mܠA�.f��3�}��Z��Z�#�-�^	W�n��G�����:l<�N��=�[����E@_��kx ����M��֟�
�JNP�Q9�`����܏�BȪ�:%��r`>��s�{������H���<����tㇽGS�ӣ�6��(�����(b�&��q)��b����=e{�[e,:�$��� �v�ݎu 
��z�X�����"s��!��Q��Vʭp+����0����)�(�|�˩ǥ<�s������r�er�R�U��9}����g��[�.��?�b%%�s޿{�ܽ{Y
��OQ���+W/�c�T�G��ׯ��LS�6&�Z�DgX�"��j�q��\!r�s�N��΃ά���܈�[��<���$���`�ɋh���43�Wp�R�ʼ���M?s��|ܹ}����O��v����Rj~G���k)�����W_}�������������_i�2���&���'�g?�Y>�����[��ؒ-$���BvG<ʎ�J�1�@�d�T��D��DC!�����.�;���~��Cy��VT��(�ˎ���'�So� ��7�?�uU�u��E	?^���Z�%LN\��@kr���#�U>'�s��)�EQu`��K�W��̲�A�&��I�R9g���Y��mYx��r��M���/��o��x��W�V���o��U�K���5J��.�4)�LN���dC�Z)'N.7�>?�����r����c�d2y=�~�o���/���kNo`ŕ$��0T�(��k�,�HV�헿'u�[������&ik��'�Vl�;�sr���S��/���R�O�ѱ1�ٯ8�,���o�+��S����~ ��(�Y�~���G$^"q��D�t���Lwӎp���Y�d��~�c�Km86���'#��"D��,����V�.�����b/D~��Ћ�e���+��
�oV8U#Wncq,\%cօ���h�]�O�z�T���<9?A�`��^�wi6��xvx���ea�TZ�RRH"��nĈ�z����־TN������t*G����>^� <4|tyQP��� ��/�] obuc�@�u�T(^��g�rq ;p�{n�s��Q!�J�U(�Y��|SA ����h�2LL�A�`D��h���k(�ǎr��D��w�J���}��	���H���\�L�ك �� @�t,�"�W�1���H�C��)��r ���BY]��)\�#�]bo޼��q�_��������Q�f���i[?^Aa�gJ��;2Y�� �L|l�������֍���'���[�ʍkg��k�ʭONI�=[�Hѽ.����k@��`(���Y�gT��S��a���������m�d�T0�6��n�ⱒ�N%0W�U��FD	B�Y�(��m�.�Y}q��LI�J�Μ�e;��rU��/>�!����W��"��O�_�(�_�b�7�����>~Y���?+�W�~U��_��(�7?����������������?/������}Q��ןIɽ]n߾^.]>/E踿��l���*g�T'����*�ڪ�����ް�3~N��-��ʼ�E)����5��5.��uO_��H
i)������e7V���o���
/+PV�)S�J�@)�XTx��E�X��Go���"���R'Q^��Y��*_��S���{/ʷ�>�������R��:P�<�cc���j+Ն.H	���Tm����$�-T����ƫ&�#c�B&���yƒR�,ǎ�%�~vK��m_��W��Ov87x��|y�x�ܻ��<}��֡trt`�� M5�-E�����c*�U�|�Hy���Y�ߖ/E�*%�ӻ�4����u�\ϱ���bye��̬��/ߔדo�\����H�z���`?D)��;���3��62_�V��J������k����N��iB��VFB�儐�Q+�l��v�����}�o,	�Ţ�Q���Rj9m��-����:��;��x 8�a>!�O��ã>;���|��3��㏄q���InQ/�g+�f��ٞ�2�����`֨�慇���v�hL��s�W�ۯ��_�m��.=� b�h�lW{,�i�fqV4Y]`��}����C�O��� �#Ӊ<eg����O��۟�H;���Сa燕h��*f���z����LL�*-��~]�е,u���`-��N�(M�Ԑ~F����������A�q�ZH_W~�uN[��At�\�q�j�z�R9���2c4 iH�N���{�[���_��dE�GG�>,ߦ����G�R�-v'�z��	t�+>�ŭ��KU!O c�
�D���Xe�~~z`w�]dj]�X�nj�¯Q���f@%�<����� �k̀���rz1��g��m����N����Μ*Ξ*�d��T����e��K���$�"��KgU�������҅�N�����f`�1d�Ӷ��۶Wb1��-������|-�������w�Pi.s��D9�t9u�t8:����
ic�GD�[Xե��O"=�����? 3�~�s�_^����D*>�a�M�)�T/#v� �\�i&T�x�VXq���������by��M��믟����A�Ϳ�+������<�Gl\>�Lf�oK1=��B�.�V���HY�ޠ�hu�K(��$��Z]2�2��󶤭�Ď��[�l޼y�\�r^��)�TN�{~M
�By�tJ����8�����:L�dR-�	���T�+�*#�:���(wQ��/ޕ�j�W���;ׄ7�O�	����is)�⒔��E����Ŕ�.f�H�xP�S�{@6́@ݩ�i/�0�*�����i�z���6�J-�-W���h��u��.���[����5�%�?\�t��X,��M2��!���#K�"�u�{�m[��GHF����ՠ�A�4懡����\�~*D|��G�.5�0e�cD�K�h���J�O�A��L��R���㆏�X��N᷐3�����G����G,���#Rl�M���_�M%,K
n�� �c�E��Ը�e@\(O(���S���Qu�G8BJ{(a(����HiȰ���r��gE�S����a�)׎ق�k�|$@�,���Fa��>0�s���+��}�T9�X9}�p9~�^�r��r�Ę��k��+(��.ׯ].G��cF(z�4X������S�V5\rv&��1�v!4@9�qǤ���5U�Mŕ�6��[�]�i@Y$=� ��3�Hd�S�JT]�'�n�L�A�� ��H�Ś�i�o�#�,��簭E�ܿx�C�b)I�!^���/?o��bo6+�[�9N�n��b����2:v���~Β])+��eaa��μ,o߾(��o�M�N�>�����˕�ʩS�j��<�ŀ4h�(��-
�Tzo�Kw�ge�&2�=򉉲E����
jWr��-��=�FM�ɟWt5��M�W%UG�����A<B�뢗��..�+og6ˋ��>��_?-��{�����?��7¯e���˿|_�����ɫ2�vN�7T��[�WI��ٳ�[$Mj85c{c�l�K�ߴ{+��ˊ�W������mM*8	c�c��xlS�rP2�(W��/�}v�|&�_�|J�ĸ�Y���s
���jy�|�ܿ�IO��/��䬷U����)Պ������HLV�X�`���ن�i[[��sS}�p�u�|����/~v����o�b�y�"��v/�GO^�����2.�����LW?z�F����JF���u���M��n�Vco�ؒP�[��
�2 ���m^Hy�6gLyD�?$��U��(j���鐜���Ⱍ�j�n�n�v��ŧ����	N���3��H�A��|��YI0��p?	Zڍ,����\�
�Q��)�@?��{�~ RE��"D��T;�'����`�XD���A�7f��C����M3�TNM�5�֠5:b��W�2K�՗-G?5�XF=��d#��ȝQ=�@e�&�ŝ�l>]��^��Ո��s{�m4b�2�#���6��,�]� 1@c	d3�_aKƜ��*�������_�)?� �嗷�ݻ�ʝ�Wʝ;Wm���RhoɼU�h�a���y����!Evqq�LO-k�c��N*-��B�B��_)33K���pnnE��t]ϫez:�.-��+�R�4))�=�{���7���p�#� E��V�uk
6jc����:C�Mj�����ֲ��]J�,5P���SR�ڣ���������ŕ� Ec~~]e���#����2'���y��6.�]��l��������6Un�Rr���su��gQR�Iʟ�G�%�@�9&����g�+���-7n\�v�+WΕK�N�N�O�˗OK�=+���;W����Oo����z�����!@�Z��/+eiY
�fWAǹ�V�s�6��A������ �]�(f(�RQ
	I�B��Z�gϠʥ���T�-�斖�
�Np����F�[X)So�N��(�|����+g�{�� ?�.O��-�_�I�>�)O�L�Ǐ^�G����ʂs����Rf���hҦ9
fw�>�-
�cp{,0H�R�	)����؎�b{���r���W]6�Ua�;
+�mO�Y*O�N�_?T>ė�C=��d�2��w���Bm�����c��:�����r��'�7���z����r���pHʑ������+)��*���<�lbe��^�_V��@�Ϗ�Z����;@�x	$Bޑ���qR��FV1����X�������7�Ŀ,X��B<�W矉[1�#d�-Y��J��0d��5P����8��Ǐ���F"4}ȶr7�GZi��R��q��'��#^�7���L������N^��^n'2m2f
������jԯ\�v�7		3��J����\� �P%|���W�1ek��==��	ǚ���������}s�	�����t����y��������WY��#<\Ν�5���I+��~f�g���bF�������~�%3���	k"��H�<ŗ�칋5�)��l-.�� ��d�W��Ri��&���%{�uTx:yM;+_MT�x��q�L����890O����jY]���Ε�������XPک��>v�P9v����ڵ���K��E0W��W������*����pO���N����i2\Q��w�����ÁK��K�>S.�;��p�ϕ�(Q3��V^_Os�|y#%w^J�������Ÿ&��+�1��l������P��`�޺�S�d��nkC���Yы���D9{�׭�_��5站��ٛ� ��零��!)�r���Z�nxU9]�p��>�y��JY�����|y�b&>�Y�C)�RLP�h�D��hnJ�X�#gF�+'O���71��]R6e��`��|c�gem�����1���'�|1��K�e^���LLPFP~Ql�Pf���	m��"�27�%J�XZޒ}K�~��>~�R�ڋ���K����/Ia�x�[N��A�����R/�o�5፛W����ݛ��{���rSn�jR�?g���CݥKb��V��{���\=y"�5����(>�:w�T9"Ypf(UaY�ɍX\ ��K�S��f�M��J�m
�,4��75�C��z��&+?1�~g����GU���>}>U<x�r�r��(�����	���8-޶���)[*�M)��ݑ#ޣ�B��M��~=�}�oްo�e)��c�������;��̖�B�/ޮ���&�M�)��{�$q�_�_�ŉǕ¹��}�����ߕ�{�r��Ge��1�)�D�����#�*nӊm\���q�Ə�R�L�sNx�����'��Ջ~C��D�	��ڎ�����O�`?2//^�͛�8��Ş`m��H;���ڿ��� |b�
[��'4�H��z���kB�GT����g��9s��78}GuNu�o8I;�7t�9���H'�k��s�;�`�*7cҧ�����A����W$��ib��вNy�G6�v�z�e7F0x��U�!J��E������8��E;�=�l���3}�q�܏��aM�8
a>�+��)��@��i�I������a���7��o�����>v�������ǆ0Q$+��j}#1�V�`�N.3C��)L�2�*S�����J��I�Vn���/�(5q3 :�����L���_�@B�p������w�EEh�O� ��PL^�#L:�3�������Ǽ��M��JE���L�� Aϡ���t�i���}�ՅrEy�YL��cKSp=
.������*�C��x$�׳��/��%W�4ă���"}��� ���{�U��6V�ڲ�[���+�\2�`E��R�8,�}tǸ���D�q�H9u����|Oz��i)�q�9WB�j֖�_��(�M�������K=O���)�(#�(��n����}m}��y˕��޳�x1�gV�^O-�zPnWz��u�|��D�eM7�^lK�U��L��·��g�%O�����vbbD��IEvFy�!!�x�������ٴ;�g���:+1O1)�*8�t�"x��MoW�y�r�t^���c�\H�UX�g��Ƿer�۬��!f{g?:�z]���؏��!�tQnᕕI�@�}�lJ��ty9�^���a)$�Œ�曷s>��Ɠ���ÛW2''�ʫ׳Ɨ�{as�� N4	;)��_�ʏ0(���&O��*�'_K�|c���
/����E���*d�8!��/v9-4�+��K�g}�K\�����c(��]f�W]oPp<|*�^Kf��;�I�P�y]�у4-����+哪_��jT2� W�:�P�J��B���}��!c5�k��r�;�2��3YS����Mf�3>`R�F�}�����v�D	�Ƹ�C��,%P	���unx�N�A	��]&dOs9üW��IA88<�<�_�R��-'����~������?��d⦷%�����L8_���d�WkQ�Q�WV���rqΪ��NKnL��֍X��b+���&���������j�|Qʵ�%�	A��[ЄW�v��+�sA��Q&�=F9����&@]�i�Rvm�������������L
7�0�g���`���!Ʉ����ŋL�5N��=z��m�;&��Z�_�|%7�d=͇��G�,Z�~��#�6�5n�vh���DoI&�t�m+z��A���o�r0?�Y�
�<n�������V�3D�����'�f�2�&����Ї�a�rK�����c�D�I�t �!�^��?�1F����ͻ�h���Ǌj���h������BI�FEl���~�C��`�D��B�e�"%�7�Q\�O�j�@���V�b���p�k
��\VLGZΜB�.0Ѱ)LZd�2ʲ�%�舣���|���qR@Є�(D�ŦK���è�'J��S'�Xϔ+/���G��pw�GP��D$ma�tp��B����{o�Lo *���[��M���~�ōu��s\M�newc�N<�y�
�tY cP�1��`C6.#��x��P̧��!������CRn�r+�R�|��!U�����rw�s�-�B��I���ZA>�C�8x;ʐ�a��v��,�o�{^���I����^��9��R9rt��KR����rLƗ�T0Hq�7�>�*��S5)��n��s�����.��ոz�,we��#/6dZf�S��yn�M���^W�ؒ2?Z._�W�5!���qd�k)�r�Z��Pn��b�+ڪ���%�����A���2�;ylBʭ|���gR�/V��U54����@-��q�2���SN�<���|��s0F�3��\�?�,�&��K��]���X�P�};�V��KM<��GR�>�B"|��P)X���|��W�>��>.�1�����BL��g��Դ�g~Ae�de���1pKye2DQO-��q��q)��O�����{M��L�<���ĸ��q��1�>�����y�ye��2���������z�B2]�,��:�̾y�&ۚ�8��������R�_�[�]Z�TA�RD��dŖ���^�R6 e�ĉ79�j�l�a��8�G�w���Eb+�K~{155-���B�/^��fW5���+X��i#�2L�>�}���P�C�r�W�9�>�-�o�.���Ԕ&�k�����(咏���m�!����j�t�h�r���ʛ�Νk���b��� ��I��GS��z����[�R�2<�|s�,K&�u��h����rMw�Glj�*�j7�2���r������ʗ�b��0�P%KV3�Puva�<y>_~��G巿�_�S��!ʵ�S�i��c*��/�& F;�5��y ����ϊ��D�Cl�B?�#���{+��3�9.��kh�ׯ^,��N����F�a˂?@t���_
�I��2m��Ya�3��ʏ��Qp�m�[>��m''[��s�:+����8=���ߊxMp�B�3�~:����Ř�EA/�NX�����(��C?*����a�c��k�?�EY�Z�ǩ���6?<��I��I�1�A'&?;�;!Ê�Wn6���6�2�m:kN#���sgO�&b�DB�40�j�t��X���f�^�MhF�b@d[���@�I�f����M �V[�	5!�lH��@rO�h��ؒx��Bȼv.����6�l{\
��$V��꫉��aF�TC׼����`�������B������F�k��2��JY�p�qn��/��U�����@�3���b��S��ԕU+/bT�Θ�]�i,r�C�V��9�AjT#G�Ud��	Oǳ���/�J��"���̒_2ؐ0ɉ���I�lKX�|�%)�3�ɓ7���7��G����dy"����2�f�,/�?P�a?_�'˪*�t��-K�d�W5���+B!�ث}Zm����*�����#�%��@�*�䧿�:���0&��`�C��b��n&C`tL�ʯ�$�(TF��������P>��� �n��n)���U)�R�_LJ�zU��<`>z:UK�~��zȗ�RT>���ޗ�<�>)��r{��U��(��eM���"�CL�����`�A�8&PJ���r{�[�d?!���'fp��!)��*��k�9)�/5�y�����g�"�?Il!ٷ_[m/�o��4pr5+�����}{��,�A��+�d���@eA7%�D�m0�0�I��NO�>?~"e�^�����<Ax��uy�v�+�[P�/;�7�я�:?����#cၺ��1���P�u\p�h26�W�n
�@�g�X�R��>E��Gn��rZb?��Ry�tZm������sؓ��b;"�(���^ųJ�6��S����V�����}��5�)���i"đf|v/�-e�Vџ��m��/�U�%��ޟ<�zA�zW��A�2�S�*Զh	��0M��o�?@�3&�.ԏ1��*I-/�W���1�M���v(�W�i��S�M��C�PE��Q�{����ʌ�l7n���`q%��U{��BIKE-*��7�J�����:�Z���S'\�!z@q)�Ѝ"0�vHO���aA�W��
��jCˑ�J�v[v�~��>��zN"�rГЉ)�H�&#Vr2̇�*.`Ud�е�l*/N*ҫI7Jm����q�'*��Ф�,@��4�o��I�J�G��C1�=�rs��v	�������H	;\�W�1��(p� ��,�ь�)Rb?�{�@e���3�8j�H>�հր���N����JSQ���8t� di�]���.s>����Z�l��,������̬y��E��{��o�/�=-�`�
<^���� Qm
�ܐs�o�:����Ux紅}B)�s���yF���[V,��o:C�bT���j�(�B�Ր�jXe5"V9�5��I��۬hn��ˮ��bkC�
�H���#ǒ�P8��nIpL搱=�A�݉c���&mK��
u���|��V��M.���N�Hn�K��X���t�(�2��^��c�Y������Dn��2|�4����#��0��	e�(#c���8x��&������(a�7wq�k�� �P��̻n+o��[�����
rN�YB��)˫k����r���؊�j�J�������D�ݖ�b/�ۋ��@A䣻�-V��m�I�g��$�sc2�v�\_v����}>,_}��<e���m%3�ڶ����j�_��b��������X�q�s{I�c��p���_�FO�
�Öx�t��R� ����K�|'��Ū�jY[��e�����֭�>?�.sV�qN$����V�O�Z.�)�}��<����}�XVWP�)���a7�o�$����C#j�j\
���
��xYT=�WN�>�7;��1�Х����L�2>7�]��\���E���'~�ª��;�5��#cGʰ���\	����\�K���:��ϕ|zA�ڭb1���݃L�2����硼1Frk^��!)�,pF��aeO���ſU Ӓ#����`���Q�cD�(�a�ɬ���o��y7�F�bB��� 7�z�NԭT����??�?o?��^�e*:ެh���s랁�(VŶ*��hl3���-d�B����k�ɐ|�m� ш�r˫#�Z���z����GV�?DAt� w��Y�(�(�|���;^�ke��`�S`��+T��� a�Z�����C��Y? �S^���3JP}eS��-�F|���L��޿�B�{��.��7��_���hJ7�����������Y)�RH�����)�E�H;os��Fd4�i�|�E�!J;�oR���&��ٔ�����*��PZ4��7:fi��;��a aS�RÖ��J�`�jR���I̉\��J��k��-ԳX�E�e�A=��+�2��m�d[��`�2J���W��?�ob#�+rb�ge�6V���7r���GG24(��q��D)�v�;����A�Ai�����
�: ����s}-N\0r-,B��i"�����Qf��z��&SϞ>������#���S
/R�)҄�~b0���%�����Η������w����Nu@J!��� ��y��������ޟ·�� Ui�^�{|�v�SU���v��e�������A�U��u=�g���6�.��'��^}��*��Հz��(���E�}�A����;n<���L�����O��z�[����Y�(L`Q`9��铙���k�I�z=�������D2yb��<ڥ�ƨ�����1��F�_�r���<�G�gˍ�}Q'�������������yo��/����WRl˚��"�p=�W�=F��BS�VBj�?v�>F��W�t��^u,���W�k��X4��t��o2o��F��2�u�2s�+�?G�t�=i�/(��p�V���aE{8�@u�8 �}μ
چ��L7�>̐{����f"üzӢ�e��#+B�S�Cb%���xw��V�GUC�#�#�_3���vf�(���&�c���SBH�J-e�@�<K�䙼��/��zt��YY��Х�p�T17JmŞzD ��!n�G��$��T↗Hip��=�*���w���o��������+����7��$/��rs��1�M�
�X�b��C\!yP2���u.�Y��Kl��Ye��U�� /�f_��Fa�՗�ź�B�gE=�B�d!kW��R�DÓ+(��Qģ�|�J'�/��fc��7��(/
�U`��"8��ie'q���S�-FZ(V(X(���d0il�+�ե���I�pme���v�W�(O����_!�Cɖ�
�dX>���Uo�`}�C�rsT�R���團����{��l�Y�ڸi
Z��4Ņd���]F)���p�2'.,n�~qbƪ&Y˚L��� �� �
�c+���r��z[�K�}��i�|9Y�g�o�䃂yX�Ha�B�b���@��_q��+�E.�X.���●7Dk�hEWe���T�I1�\�S��7/�/��U~����W���ܹs��?w��w^i��R� "@ݿϕϾ�[�꯿*��U�����|��O˥�g��##*�u�/..�8.��:�2�^_�Ū��O�	�W��'�Ue�bL$+�.d6c+�&DU�ߺOʱ��V��C[�ȱQ_����������%�}�j�S:|��N�M�yQ�ݗ�L�,ӯ�|e=6v��>\���>V��`��@��=�գ���=��.���	��PnI����)ח�j��c����M�ߕW/�˽{�!�"�g�5Mj�7$o>�ܯ���,ꗷol#3d�m+	UN{���K��c&�?���	�����6��
���g�n~���
1W�F6)Q��իK��{�@�4e�o̍2ߠ�r�ى��� �p��F'-Q"�����v|���� vܺ���M�M�����^MF`�P���N>��n�W$�z�d(��z�Ù�~4TF����@�M�aC��Z�W����bm�v���{�.&�">�c�r�GO�����N���	��(0�e�7J&��v��[�R?�磜���}��������=*���(�&�x����'R�Q����?�����<����ܯ�x�W��4��~:V	_��s��,�$y�ne+Vj=Y�����$]�����ޅR+%ү��@4C^� z���Pp�y��Q���A({^���"��k%���/�G�������xV�Xɒ���� Ϭ�w�~#����3��gʱ��e|l��.a9�[�	���(�d�+�΅�"#�	~�/֐s����P�ӭQ|��B>�7=ӥ�N(R�ޕ��u)(�ޟ����r�����|n�z�r��ίY�ڒl�d$/q<cd��<�y��u䏂5"C���D�8_��)��-�[n��Z�+��2�r��\�퐔�'�֮O>�\����Ϯ�O�^��v٧:��ܪγ_wdxD���r���_�-������R���])��ʅ��!��-��ꏻ�����r\�-�������g��Y	e�
��J�2�u�z��[�n��+�N*���/7o]-ׯ_V�=+��'�V�L^Ιf_���=+����ݷ˓GO˛�7eiaI��Gb��DAi��/*����Û(��|��O��~�'"ܺq�7��>9Q�G5{��Ϲ�O��R��|�����q����.�-L@�>����	�۬�O���BZ�f;�n��l !r������?�E�G�㪷��`ˎ��7�Y�������<E�,�'��&��͂ {��[v	�IH�"��o?�uexy�z�LP@������
�=�h���a4�v��{$�'� �Ȁ��	�$�Sa�ώ#���9͏��ex�|BS�{�#	9
�X�U�PpQ�Y!!���`����#��YFE��"���;S��'T�U�Z���3��Ӱ���@�m��R�?=��U=�b�6V�Ĭ��p�%�������ϞO��#��~�t��J�����}��l���@�8���a��r�������W�����s�؈�X�d�"��Sb�
�*,��X�E�����v���FX�ʣ��4��ec���zI��nmJ���$No@Y@Y�qy�J'-�������s��r�33�s��lI!<�x`b�lH��	�+W���]��D����L�
~���pQ�xgd���8����������'���K���c'�hk �I���([��,r����p#^ڑ��T��"|B�I�@~Pn��P�[�Qn���A��k����29�X��{^~������~[����o��!�?��������"G�Q����Vx\���r��M���]�PN�:�I�����������R(��3��ΌEQF�?��7�d��J�cb�m�۱*����bY_](�k˚m��jV8�؀�`oK��q�d�v儿z?���Lʙҡ&q��罧��P���Z���o����-�ԗRpf1��;R`ז����\�X[Rl�)mK3eyiN��^ϟ?��s���r��a�O�1C�GꙬ�?o*֔�%�\��z�8~Hm�b���?+_~yW��9����,�|�5��~�m������������*���㇏˛ׯ˂�˥�9�&��>csy��R|�XQVR�c{}e�~l����˗Η/��[~��/���.7��M�Uߑ{|9���R��__�������]y��~y;���,/(O+n;����^b�Ă��X7�1�i�a3�"�X:���6~�s`�-������T�(��e��p��|tnl�v��޹�Ti�_j��J�����_Q=O�-��������9�ɫ�ޅ��]�xDt�����-H�6.��t�����8�HС6l�+�]	��?�J��� ����zF�p�g�m������ �mE)�����j&�ȧW���|��Uk��J���3�XL=�O�`9����S5����'��RFQN'e��N��U�(C[�oH)[Y�@���9/啃�};��pv�d������OJ^P�u��SFǆ�q�jԀ��k,o��w��+W��ت�1�j�,VX@�O<aU��q��V�[o"�2C4amB(\�*qQ�8�xk���ؿ����G��'���cV�x��"�?KM��*��Ç�\��Bq��>s���Q^�G��ce耛��r�BkY��-5���F�Fˑ�C���	��=zl�9ʾ�1��<A��� .������ӻwʍ�ʩS��\�����w��x��|*R٪�h,+���S��\d�vz/j"2�s���'z�4��d�3�l����.n9��_�o�y\~����B��~���qr|	����2;��(�@�\�����d��ͫ��k�쇏����٧̞T)b�:�Q}�͆�/Տ�8Z�J�<{�d9�	����vŢ��nm���Ս�������<��.�[*Vϝ9VN+�UvyxXuɯ��6���&��O�3*�3
���r��K�j�>�s�;4>T����@���Y[�Ʒ,�7TGU�"�\�p��N�W�9��]���)�z�ݶ����T�5�r�[(������>&(Vl٦����]α}Z����������2=5%rQ�o�'�- �f�85�z��-oK�#�b�ѣ����s�}v��x`+���Α_�SX[]���/�O�G����<��Cy��Y����A)ɚ�lm�UhYyV��~�ĝ����%�/�t�S��WǍ���}������e=��!���d�-6(�U��R?�(tn_į��@'��6�=��1��O]��_������b�(��I�H;��Yk�nVlk������!���	�����Xâ�a��]���{�S�~j]�?�������oÁ^�
ޅ��6��R����2)��92����Z�3)4���u�d�#�������"�W��WB�,��w�׮(���Hɨ���8�%N�Q��Gh$_����È}���/��קc��SRl��>�dHJ�u�_.�1�~���������x�H��ݑ�i�s�Ï2Jnk����.��3���������9HJylG|Yv��?��)K�e�E�jI���2+Sn*[[+>��W���>#<t�[���XΙ]��/_�-����Uӡ��l��$��s|yE/�N�c>�6V����ȑ)i|,3�=xLr6���mƫ��DŭU��5p���V^p���/�"�M)'۬���e�:����?���"�UV�#��t�ϧN��U5�
ҵ�����g�	)�>@Yq%0g�R��v92!e����q�/勎9$�O�à���OxT�)�=s�����xX^]�
%�c��2"E��1)�j+'OKQ:�t��(���L�۷o�;�oI��&���qI�=��|�v�<y6�	���t��ZVջ��1��z��ة�U����ں�H��=��$l��UBV�V�g˨����9�9��;�cHyZ�z�%%��7��Ç/���z�-��q�+'�{*y}�#\��N� �xm�
O�������*V8WYm�>>�br�kp�	��'1�����!5�,����=�����g�x�gBs2J%]��H���`R����;ea�f��=-�3s��5��(w?�%�����s�$`%]u��(;��o�s
æ\��q%�Р<rV%bp��M^�nq��oj�@6���Ҷ��{�#���"ŉ��e���7�}����ŧ���_(�U＿U�Ǟ�%���9���Ф�kM2�)O(�+
����&8:N��M2ycǖ4�+�qdZ|<F5<����X&��ɕrI�c��rp2��ںx��b��<������~y� k�!p��?�Ƈ����(���1��o���,��{�؅��]P����M�c�ϑ�{�����
��}��?sI+�l7�7�E\�f��~�� ����4[`J"9a��z	�	m��������23�X^����2?���E�W��.n��0Q��/���W��D}��� �V�/�c3��T��������+�Y@?�]_M?g��)y���fz�m�5_�̰͘���&�*_d���K?�7��4����:��L������(cށRn�T�,>A�V��3��Մj�`���&�Ȫ�� �� f���
����&�t�e��wh��?
���.
���Z� �;v�b3Ta�d8p�6�@c�!�k�FQ$�G�Q �*Y��ָ�vE�߁��f-�
��z]~<T]�P=�G�ST���s4Xn({;3��YʭL�DV���̫��AF?A.h!w�$6v~������0*g;�N�����'���`r^J_u����W��!l^�֊��L��P\���=��(��s8V7a���`L�]��Z[_��2�vJ����l�?+�-n(�罗�~f���F�U$�L����?�c�֎X%�:����=�L�<r�=���i�/]8WN�`�h��������}��q)ħϜTǥ0����%��N�UO����0.[8��O~�u(�R��K[�\20vh��i�9w�t�x��`缔b=��-�b�B�4.Ѡ�XY��9�O���<Zn�����ջ�(o(�/�s,�|v��g�y[���	k@>�=�>gK
�Lq�Ӑ&2g��M~8���㺦�W����b;�z�����iz�.>&|L�@}�&�Y+Q2�>��Q>\�c�a����*��m0�El�2��~[�L�<��z�ʁ~�㷨��T����L�$s�棧��3|��Y��&Ŗ�Tu�e�+�5I|����k�^p?|DNT`�OSa�G�GI�w	`;���ŉ+LhX�ga�UN.�8��X�fk�-Wbs���&���9����j���{�߼����+����5Z�]�X�޹.����3�{>�@�0f"�
�����\��|m�vX�=z��ɱ�&�SR�O�<�pnJ�F����U�*�8�N�M��~Iu�k��|r��.�nW9�kH�9��������YՓ7eN|�ʜS&hW�4�L�b�q��	�|чD>�e,��z��k�@�B�V𶢧7���b�M{!OY�Ճ�#�-�%[��f�~�2Tް�V"NL�'�l�r���P��Dl�N���H���O`�$�����}M��T�1�mYXФT�%.q��Rt-KL�G=K׵2�D7�@ -�H��kV�u}F����d���L\�4�-�$BKt�M���G��N�r[�9����7�B��e��5�4�yo��I�>e7�[$�I&�ܲ�����~�^��ЂA"J�fB�w�<3Q���گ�6v'=��3��P+�:Q����Ȼ���y	�Jm-4=��Zt#�Z2퀰O�"$��-��C*0����3s�pX�:��Ǹa���p�O�X��0��J������>�G��0�N]�m�!kH~�;����e)�����a2�[^�2Xs�

�3�+�?ј�!A�a��_�`Fx��ʭY��Ϛf��R���j�4=��?�-.oH�])��c�pǷ*���4��W�qp�;)uӴ���՘"��p~-eC����{�<_�ϊ�k�W�^��&%-�[:�e�?�z�L�Y�k����D�����G#?M�y��"��p�o;��^���q5�˒��;7�_��m�K2�/G�k�eP�� ����)^%Kf.�܎j�ߖR�!�Y��r'�r�`�D��3`]�1�C��'���d38�=w��\�~�\�)^nȼ���!�� ����\KK{?�)���+v)33�Rlg�w?<�b�_LI1X��wOPT��D_U�����2������u��2��"ty��Ěc���[��s\�}.�[���yb0;���L$�Vr,���Gl��ۥP�6� p����Y��YU�\�[�k�	ا����-�-�W�P"Q��h����XV}�9&e쨔���O�K���޼�Ur��O�w>�R)����G���T��V�WVvʔ&�L�G_��/�..+�JcH������,19�Mk�3�٣{|b��;wV���OV7���9{������f�e�Rx������>M���5���K:�\�y;S67�w��I�>M4N��~�y���˭���Y)�>yC<x�^\��5(kM�$ד'N�"������N�d��k�.�MKI�r���gU�ǎO(oC��h��nl��ݹ-Y^��:}�a�W�Wun�1��	} YQ��p�&��T&����d%�>�ڍ�r�">.I�>�1�d}����z%m�
��oTe����\D���B ��c���m#�'�U@:��1gX9<�*&���F�ԁ�� :@��O��GD"}�LT9`���C�O��~9?=n�w��N��r;���W4^n����յAt���Z�� d��@�r"�17���@�D��`���#�۪o)]ד�+��{��ӯ�L�#�[�� ��hw�Ș�EZu����8�n�Qn������-��p�.W���b���g���!�\0i�H8�*��a�0��[�P%���~$���������q*M�KH!������~���`���nZX����/a�����p �lK��,#�����l\�r{H��W]\���ck4P������G����V�s*�!�i;�	�c�2��w�H9����ܶ�P~(#�IRȩ7{m��s�����-��v�?�C8B��n�X)V/�-@й3'
���<w����!����Y��Kl=���X�Bp�(3��q��1�$5XG݂����HJ�Ԍ:�)ӹpQ����'�I�u�^\\W��r;=�r��Eb��������G�Y��וY��ܘYomnh0�r˫����X�=YN��h ���$E���J)=�A'pL��29�P޾]T�*M���Qd�9���>qr�_�����Y����A�(р6!�jB
�7�3�5x��	��HI	@A�"@_��63�R�>�)�v�[_w��ک��}*;&&Q�<d�
� F�5�G~U�|˜�W�O?�q�+,u�6������C#^�G��ȫgu���yK�����$����w�e+R��Qʵ��E��E��P�Gm��T5�#�uߐ�͞q��/.���my�OA�N�z��xq�˰&��/+��4/�N��V���=}L�De��kL�#lXX�R�$��L���g�ٓIM��MʬӠnlx�G����J��L�b�+�Ú\�8��NH^�j�����0�pFn'U'�Z!b"�$wy��k�ً�������KMr&�ׂ�����\���>+wn]-�N�dn�+�4-z��c�J���1�Q��\�������e�����%���cR^'�o��xSa*���aVmy�Ҥ�Iާwoy����W[���"r y�2��v�q�:_O	�x�&��ԇ��<�#�!xs��I ��G�GUw���\�Ӈ�����Dy�s�O^�*tB���g�}@L����k�3��wD��#;V�y�9,�����o �t�J e�ȣ�Ko���+��odVT&���e�����L��K�t�X}�z�-=�V�����h��rʮA��W}�z�@�:��#9���Z�k}H���X		(�Ak�r�y3a;@?�"�Ɂ7���m9Rn5�M��b�6�%���[3X)����̦y�]���;s!4N��9	��Ō�a�]/�;��/��C!������ִ*�.����\��g�c��@����o[�e_%���`�rKc�#���)������z��np��ҩ��� �x��=��{��nI�8��o���cUvi�����Z��v}�q�P)#ńd���q�E�C&k�*A�rw��|�����p �)�^+t�ШW�N�� y�/�Ǥ��23�^^��r9�P���3g�RO��ZS��7����P��xϢ��a�C�t4�bem�g�ro?��7of\�N�>p>��0��l��7}��WS���j(F�Hp�O���#�ҮQ���O�r����:^��Xs�6�;���-�U\d\/�Y�++N�������Nc2�b��'��0�;(���W��u)�E �����N�"ٴ�!�%X�A�~�[���R��b��<y�Z�^�<�g����p�j���.jU՛���������4�z	�(0�)��_u�Uу�呎��ƫ�sR�.]<%�퐕[V�޾]S�X���E)����@E?�6�P<�{|������&]4C�?:�1XlG �x�?o���eQ�x�(�1.Y_[5NR�����r9���ge���
�䱕jT�ǈpEDȵ�t�ԏU��ٙ����Jy����垔��Wo�o?D_}�����g��2���J��ζ��
�)Y+;��C��Cl�R:~xī�(B�ʎ}��_.j3k��Mr8N������K�ڲ?���CGFʙ����ݛ��zD6�L���u�ޅ�,h��Ư35�:}�H\�|bL����0>������2���i"�*:� ��mϨ-���cVH�ܾQ.K9=&�ƕeӵ�v_��
��t�p��9�#�}>�;��[B�j�qN�ge�-������
�� � �U߳�Ğe
͔�������.H��� ��-��35t��%�y6D؀ꁞ��-A�H~��r�M����K��#(�^�?�H�#�#�����Ǧ���cՖE��^K�}��l�o��	����I;�'=9�$h�V���iWf�[�/fr-�Qƶ��U��z
�~����O�1�$��az��g�=fҦ���Qu����I$_�rK�O��g�v�oѼ-�X�a�2-t?#�����M4�G���-���d��TL���o6гrkZ��$��FԦ��-B��;6��Ii@�E�Uc� �>"����v����HB�,+�u!��@uK�A�{��:q��^���.Y� y��Un����-��H�Et
�J����Z/����iX��*��F*�Qn�/�{!7��7qlB��W�o;�,c�<y�F3�9u:�V�zh�����hZ��|PJSU4}�����U]�����ūY�&���5��9*%o�8���ߕ������J�+^�]�6u>�>"�&�Z��&:�m�,����ثȀ�>H*W�n�\�@)S�O+sc�7 �+r[Z�Tg<��_s��x��7e�DP^|r�FmVf�U���Ƹ���"<�������4J��P�QH}��&(�N?yZY��O>��r��<y:)y/x�-��rSg���ʋ�ҬC���'�6?�2W�u��QBh%C?�#�Tٚ��>�C�g��_��Y��Z*�4�y�򍷮lnhr���:p�Oi�g¾!Eis����5Y���x�R]ZP{{�j�{��P�7)(����l���Ό�+�0﷥���GO9��j��C�Q�/��r���gOg�TN�{?�(�N�ׯس��"|P�+����5��>���E��ѦB�f�]�6����U��V
��by�	W˳�s��}nj{�v��ۢVָ�a[q���'8��L�v�R9�AnY�$�e��'m�S��t�2�y�|���j���j"ǖ'^��Ȥ�qz�W�&_Y�gk�F�n^��zxL����Y�m������v�C˙���_>�dLA	<<.w���/^Qȩ��4ϭz{ȼ&����HùU^��tk�9����o�����<��.R�X�e��B*VOX��q��ky��GlQ�?�T:�t#wd�3r%��hU��xm0�"�8�L>xe����)���jbN�n�q�~��[�U��#���P��}�}F�n#���_�.$~*�u0�[q-h4t@�'U��_��ŧC��a��(�����a �����&6��~�t��*����^�[Vny��~Ώn�[B҉B����	���*��±%�
[M1���?�(@e��ܲ�ܛ�ML:`	I���-���̓�߯�*R�bƏ��ţ�ˏ<S}��ȷ�!ʭD�^2:C+�lK��yu@��oD#�k3��J!Y�d�ו��7�}��AE遾���^i&G�W�\5�R�&[>*[X�`ʶ�)�_�(�@���!yo�t�Ҳs����F7hu�\��`���^F^ٲJ���ty,刳m��g4`���(*s*��G��2I� A���AtiyIy]�G �����'��|�,��� 7]�4�(�|�-xxX�>�E)�3�����>�ʉu��	�Z�ZY4��s�AvL:��˯��t<(��#��פد��8�l~Q��Z��;���F�]X-��,��Oߔ�_J~�R���xu��m�/�����M��$/��k��#���cu=����Rb��6�H6�ĉs⅛�8T��C��z*��W�WES%\�G�%��2������0�n�	��nt=�J�3(7�����X��G� [&ܚ���D�#�Xee�S�׬�Q��!|%��.u���U_�$�N=���r[��V��uM6�����nЀ�n�ȃ���ج0#{��uN�+�zF��
���?�U�֎ʉ�è�E�2�&[8��)��_?,_��ܿ����$��
o2FF�d�!���d����U�+�u+�!AR��v�A�捏�6�I��Ch�����7oV���H�}Y�W��^LY���Y�����)��'���g�ͅ���*AA��g�Q�z�$�`���g`[�d��䖲}��iYY^�2:^8!�����J��1���$�D�~����E6�B'�(�["�[6��j+[���?yQ�f��Oa�'��,�nC'i;L�����d���ִ8�JTmV
�,��W�!�1o�`R��%�)S!��@���G�f�q�X��q��P�Ar���~ס��YA�b��Y�_*Sof�^_��ۉ���H�í�j��>�
D���"��*�Ӑ�˶a.f�m�W����x�	z��H�C\��Zw<�Z�V�o�9Y��$�h�M;m���?qI?U�~�6x��2�0A�a<^6��#Qn���rˤ6�[NK0Q�`��ẽ�2��\�c���L44:��ՙR��Dsu�b��C.q���=��_��B\=q(�<�$+�mU:t�X�=2��LK=���(�P��` O��/�9�Z�����'�WZ�H9ބ����HQ���`Z�� y�t"��n]w��
�'𴓸���Q<�o��򱘯�D���+S(�3K��hCu��[�i������у��?M~lGd���joJI�I�W) y���9��Y3��PƗ������)���v苆1y#�NUάF�	W4`�t�����mF���J���L}+H��x5Ŷ����NIn(9+��m/�bÎ�̹f�2��N?ʅ6v��p��B���
����ry+~�Æ9�ߤ�ɩ��JJ���omN�~99�/��>���`A��t�|hCH�di;b��6�-�"M~��.I.����'k�י#��� ~�O�U��K��K���ыK6^H��o�{'ő�ZVm�1��)����1��{�sl�	U)px���� ��Q90�����Pnc���Q`p&��ϳ�o4�މ)��Ϧ�+�S�v��˾=>JY�R�$rvn���=�`�:��5�$�ʿ�HP��n�?�®:�
:�/�mJ9V]��@�[�ԖUlu��L�T�'��d�<|8Y�����r�CL>&��V[d�b�A�!}�+���~=3��dG��?�T^X��83�Z楴�-����iMp^M.�'�ޖ��&ˣ'��hefnъ-���N͝&Ģ[b��x�}D����&Y�7�:O�<�b�rL8A�@2ᣞ/�\�D��L��"{��A��H�G�\����啔�:W�9�6�ce��P٤��g3���8�Ř�#+����Q�p�ֳ�lE��.
Y�F��yA�޾�^���/��6�ޖ@�P��լд�.�V#��e�FP�I5� ��� ����r���G΍�c>�a4��ZO��tܞ�/xE��#g�����-5����p"!��DƳ��c�ڊ��������ó0��<\D����c�|�o�|{�h�_ 9�Ǭ�}�۷u��h{�Y�+ri�[�ѦnZ��o�{j�H5�X�7(:ć�u7a_}�-��xl���Pn�&`�Q_�����7i	�ϱrr�N�r�����v�7���?�t��W�����Z1e�()q�:�-uV�6��7�)�whd���{��F�����U�d��/�}e|��H�*;�T��O(拊_~D�ݦx�	�4؇F����f��#7$AtL�|L~TL2_?��;�.�6�N��,}ok�����< !��K��kWN���.�˗Ζ�gN���Y�T��S����A�
f��F|E	��z�Z��`[�*�� �G��ߒL��Li�(k>_rӊ�w?<-��Ҁ7-�dѝ7���Y6Vo���!��`x�]�V��n��J�����'�̘x�rK�Hm:���8螽�Y��#���ɖ,.��ë�X���+>(�\V)yu��[�m�m-Ы�$�}%��E��u^��|p�)t��-v:Xݫ[�D ܑ%]'3Y�d0a�$�*�*ٯ��2^�s�ɞ0��g@f��j�=x����l9�#���ϯ�Y��3B���2������Nnט(�VH��s���&+�V��\y�OJ��{����G�zEF�o�	�����\��0�_L4@h�;Ccs��2`����U�꣎NMx�:�)�Q��� -i��3� Ԣ�A4��eu�>�
����R8=������IYDy�4�[ď�a�#��Q��y����|TFz�?�)?ʫ���A��:�
>�\V��˞N���o����6�U+�P������J���O�(ǏOh�9�W�^�P���,�&�,˝�d�^��;7�(\�2�[���%�'�t}ܔ���q�/��y������KM�c�gI;eӐ�n%��E�����n�O�=D��b�|�	�&��'_�6ʑ�����>c��)}����Yh%��E�M�q��!��?5�b����/c5�	+��1�{��E��䑳S��)�Ȉ)4�\��3F�_�<�[��$⹶�t��
�k2}�����Mq�!�c_9>1�[?�u���䔫��x��6É!��E�����B��[9���K�gt#��e���k-D?!7GP͛0ܡc4�>u���`���l�>[��UDJ���τ/���[]�D�Dg��7
L��o%E/ �-QH�|q��A�Y�M�͙'��S�ʏ�)�ÇY�б����6�h��w雭�)]�x����@��3�@K��cz�d�Q{Eg�[�O�8R��Ď�%3&�O�t�#ޝ/�m��'/N�i�1��ޚQO9��Lv�WE{�?:R�]<]�~r�|��;Rn�?��&7�!���hd��+�Å"H��cjF��CBbdc�S|[�r�HW (�"$w��`��v)��H�H��!8��Ԋ-���ܒye��}[��(HB�r�D�^3���Rv(t��z�f*�J��� ����46���/'��h�pD)G�\(�.����:�#
�V�΋z҇^6N���+���c�Ʋ��k�>�KV^�c� ^�(P>L�η���7�=7x=z-�ly��C�Y�!��A�����I�L�"V����G'�f��S`�T*>Nt�4H�
�em�U)�O��⑌"�
G��z�Ζ���TnF����U>������ZW�S>�4vL��i:A�/��H����W�d6�d�j��2�tM�`Tg9�3�h��M���4���~"��0#�<،��Y��R`8��?���c�y�BlE3! �QDL�q��Z;�n��:A��c��� �+/V����*%�Ɍ?�S>X��,��������U����t��(+����>2;�@e 呕M�D�2�>��\�<�)*s�Ao3a��}ݲ�j��­��e�#�����2��\h���I񗲩���~d�u��K<�}�&̪��g�6�T�!]����{wh����{c�c��[L�Eӊm��W��V��t�W���>��I���E�s����C��Ϝz�5&��#�"������H}~��qCհ��C�h]�P��ovv�����~ｦ^���$�Zw���GA�w ?��x���Wi@f�����r龝����r��D�������哛�|��X�qx�U�f\tdJR�)�Pn�K�B�~n�UnMs�௅FD��|Z�eg*�Q��S��\w�>pv<x��Q�佼��QO�O�[��^�'Ϧˬ���R�9I��o��Nպ�7I*[�8@�a���[�#ޖP�����(���si�A�e!�+�[�G+ˍަ��ת܆��q��Ϭ��s�\��ֵT'IߡS���xr���'��\��D�~�<%�z��7�bz�VnG��Kgʧ�\)���n������"BQuƂKGE�!I�Ӭ�"�FH� ��Y��T����:>!B�C��r;,e�T���5+�
T�a%��[��4 �[^�+���¯�m�'��Y����*m���Ox�)�����k*���G�ʙ�ܧ~�\�|�gv޸v��:q�p$y�F
�皾[�(f�n�����>j��F-�~�z+?�.���T�����9��^ϗ'O�˽�j�29%`vfU������ �[���)�j���������P���Ϧ[H���?�k���#�>Kơ��� N�Ft��ЄGm���s��.�j�%Ȑ(���r�M��&^:az��l1鬜�x�^8LG!\�Fd�?��B���v�7;*�EǄ>�F�v��!�� ��dF�������V��<�zDv�"�]p'O�@?���e8?G�A�~�o]��ĕYYHX���@����
�i؉p�ԺV�xN��#͖����� iJyU_XOypyQGh#��1d�Vʕ!V4CI��T��,�����Ȫs��E�~S���'���H&�]���'L�ǀH9�5���;�ߊ�D��>zSJ0]�c��t �Q^�N�1٢��~�]�[٭�8K�[�X����K��1�9��ñ�>��&�hW��沀?�T��r�:d�؇p!�Pn�}�&��WYŗ���}1q��3�3�����y77� ��t��.dz�P�\Vo���#�3O-�4^� t�ƥr��)�*��{b�H9����R��Q2U6䵋���]h��H*����?����<HZU�8ș�A}Bǐ�Z��ˋI��x��E��J٪��nH
���͝�cN��S|��d��ϪV}�it-�s���Z��C��$)������ܡ�1f��LΨ��Un�'d`	��Lm��6}"�Es�r�v�0���G��������(��Qn�����S����1�lYy��g��@v��DTb�9nf��=���
m�`]�T��ǌčZl?KF�@�
 ���+
J�31i9N�C��tp�ڤ�2:����B@����Q|����ˑ:��c���8��@^��*��Vp!zf	�|6c~l�k�=A�00
���_�`�W:o�2�g��.eie����ڟ}�33Keqa]��[ �_0�Z%�������	�F�����t;��a:A��Ɇ�7��.]Jh햞�V4�p���0`>Ư5*D����I�M��'流a�-ݭ<�_\��rw8h�"i��A�dBB��L�=���rZA eg2�Ս� M����T�i7��Q.�Z���[��g��xE]v����B��y�1y$�AP��T�U����[7Ґ����+�s��)��a�&���2�g�� �vKރ�Pq!�2Ph����Xv�W�ZH��WOa�=���r��U�0ee%VA���m>��H�u�������I}���,���c�XUe��S*m���m���M�Jc�)7��� @��&����y���f!W��/B����������E)<�K�/m.�G�r���}���s"'��.sa�>�7e\���I�CJr�n��N�g�)��{��~`��M*-4lk3&C�)D�+�x�x��|le�`�m��w���<3;~��@�r�rk�L�B6�Жu�o�[f�����k�m'
��|[a�^�xJ{h��L׺W���2�k����<"� �-��d�	]%`}���AS|�~Śi��`���X�Mz��iQN��8|Di�������KU�qpT��&�O��8��lx��s�wl�V�*''����g�����GQt�50O�� ̴�F��]L0��~�eE�f�lBYH��(�*@ŷr�s*�Ӈ0{���а#��B�
���T4���y������P�	IUD���~pfR(�4V^s�!����f�8���X��
I+�k@f�I��vљsJaVv�1~��]�ա���#�e
�xpLy�1���f�c��%)IףR�����`3�r�a@%XqO�x�s����Elp�Si�Ҭ���Q��A�t ��x�؃vu���5���{�c�Y����x�~~ĞPUhQj��.�g�)�鑎�ob��{�쀐�Q��o��W�xe�p����a���k���:�0�=n�z����À�Nc@���/�.@�"��r�2��OV:	x��h�mQ|������!�~�iƯ��E<�06�}*������?�L�?M>L7	F8��
+�K�:�1}�#��j݈���cd�鹞�D��y�LM�y	FYv8����w���&��լ��JS�B�[yCiS��W+OJ�mD��$�mZ�C�W���}��62!L�W�<��e̘�!�(#OdG�|k�:Ș�f���S��ծ]g�݅�2{?�����K�O�Fp&cV�~�a��K��2��K�Vl����͛�C�#.�,x��3H
�H,�63=`��#��|���E9�[ď>*��:޽�k����#�^N��89�rf6ζ�D!�����VnS�Ʌ~B�n;�C��J�m$]�uIa��-�훶MیDF�׻J
C<�@�r�%��m�g9ІGJ� ��g$!у���  �	Ш�đ;�*ʝ:᱆tЩ���6&���K� �\賧�~w�4 7&2@F� �a �T0'�&�D��	�t`������=�ߓhƠQ�v&�?�!F�U�I��W��1Sې��yv̸���7��{��&Gl*h%O�1�1v�+)9�S샽�?���84Ϛv�
���n|����'�W��r�ba�������\ Ձ�$~ �2v���VC��n�-�%��Cq;�4fb���f���	��_�<�`�N�����m�}TY��n�(��C1����
m�T$:�[�ǃ��S�C����<ʴ�,�t�@�N5�*��ď0ͣ~���X�s�կ?��W��4�����i����:���J!��
}
��c����u/f�q:�5m�VeAaR1�J���������}O�ro"�l�eE���e!�`��\�2<:Z��h��y��m[�zP�A�7��Ko��o�7��Ȣ
��#/��}k �iW���<wP�b�욷 M9�
�9�~������@�Qk�$�'��%^(Y��8�SD��hL�_)K|8��ĹO�/ּ9'�z!�>�u�)ܷ`*"�X\�:V�_D��	
�k[�x���^f�8fV��ꅲ��$'�����e�=H��r$�ț���#��|���h�~4T>l�@&��dJfw@xC�=��@&ڃ������L9M����m��蘼a����f
=։%��Қd���A��ׇ�4mB�:4T�xu���M�,h+�j�Ld�?�q3�������+����!	���ZE� y�D~�W��?��� ��W&G��F�|@v���*��:��hfv�_,���������?��9���n}�q
���q�l�k���C&j+�J'������D˰
p��#�u��#����T#�@��{�4 �~n�Q���*H芏~e��e�;�`*PIӊ�N�O �K��PeCP�#/!�
m�#{�}�Q��=�v�N�[�)��2���/v���/^Qr�%�����IY:n��	G���y��R�z�:"ӫ�B��E±7oc�pc��ښ/��G͊
u�o�e.��V��An(��*8���8a���EZ�6���o!�)��Ć���1�8��*ݪȊ�ȃ�w��pX�f�dV���V��	i^��J��b��P��E����S���t||��͑��N�v<�O�׏��O�1`$%��bEi� ��Y��c<V4_OϔW�6!�p�#W��A�H~�o�k�N�!k�)��_�Cx�GB��:u=�i�\A��^���z�.�����K��h�W���R��8�7��)0x�?��"M��]耆��P�1;a�xP���oV���W�N�d r�y;~�]7?���䢫Q�I�<�C
�)��=��ڑ���?*�)XD���5\�6C�̿�#ak�Jl]p�NX�;��<uy�< �A�k���֝?,�|����[�����y�f�|1�s�A3ȓ�X�b�1
#���D��]��������⧼�~])4/B��J���ٹE��r+��s~f��:�2Hv蛤��o	E�p���z ����&� |?d�2"l�֕�O���i�З=�ƂQ�Z>����n݇��࿏��V���GZ�AyT7:�x��(G�֕�����������*�ڏW���'C'���`�[ĉ�[�����u��$�"�~l�(0B�~.��1[a�WA4�6��t���F0�4�@܈��:��'l�(Z5^�MX�/Q0c�C*�Rv~��Q(=	���~�~��3���T��b ���q�:�ş������L7��������{̸�E�*�2}BH>[������ቯ��x���7hfj�o��}�!���{`�1�[���.^8�w^�$�_�G�q�6
�<{�������3�zfO��Ig�=��u�p]��q��Yr�%�xA*i��!<�Gٲ �.�V76��*�,�7�se��L���(�g��*ul٣M�d�[��<S�Pl{�퐘�կ᭖kG��C��]֌	�1�e�;q�$����5�耮˔k��N�Q��Y�o�㪰&.�V���	�����j !�Zf�<p�3n(�9�.��'d�`*L�6M��d´{�)��CC�̛U2j��\|��"i�@���jB*��";tb?l���Zv@!��#�x�o��'7�V葒h(���?�H��C�@MWi�~D����h�_�z��S?rs��L��xFn]$@��v�#p��� A�����\rp� b���b���܈ā�sq��oZ٢s���JNܖ=�#"�$���]�
yy�cA��/d!/�k@��!�*�����p}���3�37�����;P<��A��1 R����֝t�
(u��f�"�m�a'�K��#P5��g��s�p˰=�[ǿN�mwĞ��G��h!�lΨ��'X�{C�������s�6v �k~�7_�p���.�x�N���ԕ>����Y�m�"݊��2�4Ѝ/��W��F(�o\��M(���&·��igW�{��b_�AVQ��M/i�$���GP�
��L�(��@j���Z��*2^�8c���0]�1~��	m���>Bܫ|�Y�L�'�9��w��	ɷ�^i��������a��=����c�]v�C�x4Q�F��N���An�A^_�
�M/���%[E�uz4]���v���e�#w��(��L %��׉�~�[}#��'.E�2���D
����=���H�EI��A�ss�2��s�H]��2;���Q`�n��٭۠#)<�xo�Ϳ���ѳ�B�A��I�����_�'P���%���K�}q�x�zV���u��'@���bX��	ٚ�y��H_q���!} ����Wnl��|P6>ƞ�#���c�ܙ�qC��_�̬3�k02�Vda�l��Kt�#.4�I�+FE����!����(L�szݠN�)�Tp���g$�
' kW�V�������]>K�B��D��9�����b��a�OP�?�7h��2���u�O�����t�?B���s��h�\3뛸^N��rn1Z�_mNH��lV$�$��d���f��pB@����!�����Q8D�n�� ��pu$/-8��8g��({o�	--��I/��C�P�N̕�E�0�?�:�]�4��J��t��5���_~j<0�3=�C�Q7"o]�B��������@����UN{C$��|4Q��䎼:n$ߔ���%��;��jY�cdx�SP�i5�p2˱[�a��k1fxv�r�@�L�t(��iZ�I4$]��1<����^��G�[��-��'���U�0W�d�~���_�T{}����?	�Ͽ�}�'@�.����O�L&�� ���1�`��<R��6�)|��ee����p��Hp�ճCLӈ2k&��U?�ט�D�
3�i�!`Mۧ|l��rK%7ۭz�����_��Ȫ�T�>{��*�=���ϰ������z�i�w?���-=E4�Ŭ��O����DX=�C2�,�8L��&�߲s¢�@Hچ��865t%|��������Z.��� ʃ��ԋ��Y���_�?�m�>���J��*���p���r�ır��))����?F����(EX�X`x�N�g�L�؂zn���	ނ�r�t��[f�)���3��`*]ū�tWn����|Q��'H X����d�4�~$J�tg���@���"t+����lPj�Yȳ*�,^�4*�-���nH܈}7b(|#��@���:]�I��z���}}�f�ϟ�v�����uͬi��4^��J2ͤ���g���f'��=cT0�{�{�*P^����Q�� {�2��Ϙ{$�Q���Cv�A�D�^���:����1��N-��-�8�%$��D�l�?ɶ+�;��F�PN����#�?x��6 ~,O"U��Ȭ�g_���-�a#ݱm`��1��4�U�ڗ�!�M�i�@��)J���0��v黿��tm�/�?}����Q�p�Q �tM������$�<a��Ĭ~u�z찇1��>Ǜ�|ޣ�3/�$����c�̚��`N��M}p����K�qL��0���?LV�}��n׭���l���7��8��?=����?�����C�����gʃ2��7���7.�P�������q�J��_*�Rjgf�J|Nc���r�5W�.�s����)��vs��	9֛�4l�he����Lo�I��:��<"�&���˂���$�xK:��4T���mK�T�h�&/��\""s�O�-
!��@�C�A������\���6D!:��t@;� J$��$��ӷr;z������(�^�e[T� &�d"�c��",|3��S�f(h5���:tޣ�*���N�y�]�xѹU:�-A?�/g'�gT
H6�O�:���b�m���j)RY�D�?���c�7OB��p������O��
�O���=�����6
F/(�&L�9f��M8|Y�-'#�оz5]^
��~~�� �G6�[�-�i
I_�J���'^����<x���7����C����a�\W{����	��w��O��{0��2�����|Gy:��h�h��MP�aĥ�����Pi����@3��]���I��g������� _�2I{��g{��ˮ�����
��>��õ��G�
�64����?�2�#4剿]2��a�w{��!����G0a���3�-}��y�!m�� !#R�h�8�ôȟ������$ϲL+�7�q�N?�H�tp�߰��	{F�C|6<���a%�r.����v��X9e\"�
{`5V�q�c�p��C|��J)p���Ǌ��<�"��+6J��y�+�+��e�ֈ�w� �a5�������Pp�o⛔�Tl�w���l[)�)�ΐ��$=�J'J��^�[�����[����k�i(�Tn��^e��&iTn�P�R?���K��ل(�C�w�ق�����حOb�/A�@YS�x�|�G�qM�Q0��^�Rf�]�r{\���-ᢔ���c!5=��sx�=3����)�(|� ���S�t���HH�
EJ�B����o��#�U��$dZ�R��Y��|��!��vnG#�o������ȳ�p�*@/���%d(��͆���!��5�<��?��J����wY��MU^�2�T��So��N�~S���|����$0c�w*�A�4ܤ��$��z�@��G�e���L�3�ԑ�gAH�}6���x�����}�r�@-�A�r��6����N}������W:}�ߓ�> ���t�4	�qr^��ۚ��>VP�n��_Ҭ%��I׿��Cf��ƱI?�*a���~]�w��N����2��|)|D᧋�f8��o�s��f��ڏ�8j;�Ú>���#	{�o�~����k�ۭ���ډ@��Ր_.6D�ý
ؤ!�K�8�0mHԱ���v�2ރVn��:�q�5�`Z���P��`:�0�c��+N���`Nm�|�cW6o���&F"z��D��[��T���-N��&�Pf9S��-\��ւ���^O��
.J1{|���×k,{�vݗp�����[N��9?�s �//�����s+�*c��-	ΐ��1t!�=�	�CD���*�}EX���m(_FVo�NX����[��q3;�%��fI���dw{c[��[�r�=�J��`�ƨ�i'|P����mz�K��q�T1�;���zHg[�ۣ����=���rĈX�D�D�P(�0��VBN̂��̨#	���L� ��VyV�ʆL��분��o�ū�t��ܫ���R+�̫�d^��;o�r���]P!1	���qp'F�.d�X>�8�_qE]�����tRf
�l[>�0�	V�ي_�7�͚���en+({l9��F�z*nW�NI���Y�b����R*��(��%�Y��Nv�B댇Y���1q��[{����l�z�a0��{7~?4u*�ϻ�ܸ� M�6�vө{�h���z�O��W���A%D���ǃ��&?��i�M/��)lQ�]���O���������DM���Ё�(�+��:�u�tq7�~�����������ï�h�S]���^9����4�|hHS�Z?����O���<+��0�B�vAPL��;d�p���� �w�P�+�2����f��D���=c�]�c
�VŖ�.Ծ��ϸQ��P�f+�[{G��=�`���ï�* ��J鑢�cT^����P���U6��!���QL�OVcv�R!�;g�J�Ì��֟����ƾ�͎��X�ek������Ū-
��R���t�ZYY�5�C��#嶫�fmH���A|�CX���q�G({��7e�!�$��d���ն^�E���%Ft����}�L�l�&��-I��W���[�ZQ#B��_y�	bb�GoB\�~���>���SO��e}٭�(ǎ���'&�����6�p�snC~I��L��u�R�u�����D��S���U����9�ʭ��;'�4�옼$�F�>�V����6�ä�ʦ�(��_�*����6�z��Y�3��i������q�l隗Prkŭ��B�O.��DxI~@�w�I�pT��A���+#3�}j̛eF3ҩ�������b�0��tĕ���W���o�QYP�T!���<���|5�LU�
�`�]C�&�W��=�K��	u=����7<�p tx���>�x�q�CJLX�	�`Չ�,�v��������D�@�f�!`��K��&��	���Ԑt��L��'�[>�������P�վ�K�>�7N�=�#�eهU��`�w��`�]�j
�j�oo���E�B�/ծ�P��׉��LK/���W�v'}�<^T�qON��������>?|�/�6��(m���n<}��H�y�v3e�d��8Q*�-T7�4cF� p~S�����oh�O��o±�3C*�-��n�ۯ�ل塓�1�%H�fȆqQ&�"RRϡAbFIdŊ�&�)�纷�g�ǆ���mH�d!F�익"��a��k�W����5VgQR�zyմ�|�sޡ�9����UZ)�U��
4=�i�غ|1��0�� ��ќ�\u��� �m���H�EP����eG�D&l���V����^A3h�� �c����Qn�F���q��j����m�3A�p��	[��ټC��"}cggC概o�юr{���Pn� ��L�(+�tP����#Y �Nd0�
:x�;t��� `?*�!GO!xE(7>q̇l"(�ڠ���|�hŏ��"_�iY)���u��2a�N�k��	�.�'>(;�����3��C��W�t��V.#����DE=H��+��~��
'�Ȥ{�%�l1)�_W���iVk9��;�'��N�NΕ�7env�,.�Y0����}/u;��ʁ�M�)q�tʲtM 3�0���?�!0����n�U��.��+�H���u�3?�����[���sE����v���^�K��<�����v�^lt�D�c�f��DfH]f�|�W�(�H���cRܲ���(T�M����
&$�[����,�]v��"��)�p@5+�~.�.K��;?�e������zK�k� �o T1Wz���+��\ ���t�� �������8�}�~�:a��0:�i26%!C�k!ND?M�>h�%�
+\<��o��&-a�ٲu�M�����笵�	�A�!{�L84�<�`�����p��x�5��_�3��l�ۑb��Vf��r�:ʮ���kC�QY+�k�C��%5��[[�}�~Nz|D��^|8ƾ[a�F�?�2�Ӣ�b��./3.n�m&+��w/�-��${��&�L���0���Qt��A���D/�`�J��3^�.�F�N��(�k�� �Uo�4��c"���)�Q.��;�9�9@��fK#�&o�A3!f�#�W�:/֔�BXhUz&#{���EA�nʠ��!:�QH�����C>-��YNK`��r�Ҩ��`RP�6�*���QRU���ps��!+<t$ �VF�s��rMs.D�J(�aE�5����@aǫ���:��=�!*�$�˜��� /1[4ɴ��BE�� �>U��3ܜ������CnС�PhF�n��5��VVd ���T����!��
m�s�}ʂä�`lM�}Y�S^�����"H�}9�y�l�_.���RG�N�3g�[�*b�&~�"a�q(�!������Y��A��h���Kԙ~�@5w�����k��n��=$V�	c?�(�Ο��_�@�M\�Y�tÓ{���� ҡ���	X� ��:�#2[��N���u�ړ�4#y��<���TУ�*�Vɿ�1Aʤ�K��{��;�v
�W��f� �w>�^�"������XшN?&ҕ�����tFcn��!;�4k�X��8��w0�z f���`�Q ����'&�oP�ڴ�����v�����R_L���w�ͳb���#+�|%+� �F�VD���I�|������֭+�I�4��ëB�Z2�D�MCD��2�?xe�J�x�P����*�<��ʺ
�XIS�e,vb��du~p2/�?�S��on�JD�[6��]���3QV�8z���0Q`�*-�Pf��K67V�)ss]��Z�q<O��m�E��N|̰3r�~,��\��*�H/�����>-���(����w��RR��"��#�J�BL㤕��1�ת<��Z,"a�)~0��t�W*��JX�
�6ܨ��S���Z׳	��	%� �4΋޶d���Y�[�u����x��]�!'�����Vn��-޲G}DN�bv������^<��r���[�;XNN)gN�r���!� �|OC��f4�(19��Ǘk�l��v3�Lb�9��%�@�"H0�6�li9����e�*x�
�.?�L`�� ˴(���B<�W�P��n����<��@ބ�e{���v��6���?�?����@F��1@)9�GJS��#vd�ՇEŎ���[�r���ۙ��7Rr�S�]�bKV��Nǡ6��_�(ɑwJ�B9�b���I����Te9�!U�X��[����D�\��3��� 7���.ؽ'~�} �8�l��K����	g��ʵ��FK��B��:�v�:)�@����{�ec��lf[��iS=�rd�s1���e������`�R�{�c-K�)��j���|mį��<�O�����#�^��0.wh�8��̆�2 �Ս#�e��SPe�8��� ����Mq{�1�r��� ��MW�լϤR�"�{A~5OFP�F,� ��S��12az��@�~�O���03^e��� �xnɯ���-�B��K�u��_�h�9�����%M������w�`>��{���Ä".2�dVpy����+͑7�(��3+��C�E�e�6�*����p�nRL�qd�vy��-���V��"[V����ܗX�E��6�"���V�r�Z�3����\(k*+n��4q`C�2���9&f$��'yT+�Gˈ��IO(F a��"��!AyT�6�=�KA��e;|99��r���C\O`DK��5�Ɗ��NuoM0�9��tb�v���Z�=�\��*�<��
��b��(2'nM�x*�P��c���0'�M2&z��CA��F��ҊF��/J�D��t�J���?�6R�l�0d���jC��N8�7��<#�B��l��d��]m�4VB~թJ��x�ZFu��?0!T�T�!$mh�?�����ʇrd��k�(�ӛ� W4C]ZҬta���ƌtn^���23��j�lEXfՖW:t0�*PG�!G'N�t�2Z?�d�O�Q6��\��w�23d<���ĳb����P�D�D�� C��Є�HpYd~?��q��Is�W���ޟ���oԑ�����r��pM�|�Q���q�W����@�i�����B�mc����3�	�EH9��J��O��&t��#b��C=����K�0;e���ynH{�N���i��� Ni7�=��速:�-[̏�����OoP��B�E��R�A�������&C�+�J��v�Q���� F�<�w�
���q���dE]u�1�<ZA�5�:����������?����:lb��3��:�� �xB�cdbф�Š؎P��Ve�U\�[�$��ZM�\���6�k��x�[���$�/��`�+��[�Jn�\�m��k��<.V��c#c"Ұ��v	7�n]�z��o�6�S
0c� AY����|�>d��Yȓ4�?��y��f��$	+��4Lۅ��ϫ�a��"v:zn0hb'{�[Q��ݐ�ȿ?�K���U���U:a���r���snϟ9U��&#e���.+����D"dE�f2�,a�"��R;C�Wn- \�dzR�0��@�	�V���[��i�@�	 %��j�`��vs��#ݡ�-���r0�Mȣ��k9�"���i4XW�	�RK��L:Z�i���/>y&LU�c_+4�g�q�u�Ѧܔ��	7<2�,�xe��=Y�]��������m<=;�d�vnnUJo�'ZS^�����V���;��Ƚb���)�����&X���o�q����N� Y�����]$k��v�}���
p0�x�:�ڍ{-�j��rÄ���8�G���%�ne��?+F�9�O#��?��^��i�>cZn�ว��W��?��S����P���C��K����[�캷���>p^:,5�� �t�,�Y��S�/n-��p7(���t���t��*c��" ~�	o�9��I���!�4������q�J.0[�SV�C4N���S��U!Pp�~+4�G -
;P�l!n� �x�CH+��[]`YD�p�1(Vh�:�1S�B��=E?a�W��.2VŖ-�~ ��b���"G����f���2&Z�e��:�5I܇�b�oX��y�9��G_��R���:0��2
�?���e��zO��x��<�M ��°/�*nu���������Y�
!�*���z`������F�"Q�[�Ե��[�o�<�nʢ�-�	�ӏS5�m��+�[qC��	Vn����8-AH��1�����h78�1C1��VHM&�����r+:FV��	E��Z����oN�&f��t��>q��naw~;�<����2�R��*D�.��
��6�m(��:��B��\W#��k�M���+{�6�@}4ɺhlv�,>��X�>�U5`��\�������
d3�PJ�۷�ezz�W�~=�[ȸ�7��ScW�gf̫!���\�P�o����h d<DE��]��MJJ��w@����ϩ��Ǯm (�(����t���Ww>}�4����j�{���{Gr{�x������_�́e1��Ǻ
�u��>�f=@z`X��*
���

��a�9�uV�N"�<h$�mv��[����q�c�!�OoO�xt={���{ �=*�
}~���S�M�GB_\��8��/�Py������"�}�wm h�	��u1�r��7�3�� ��>֘a9�'d�>ȱR�O�c������lY�����~�H:![L'' L�y���S�fӲjpYھ2uCL0��x�NcQlUD�Eь�	r�ي����FP�k�T���^�;�|4�6=[L��8���+��!ކ�S���<J8�I��ݝQ�@���=��y��)w+B؅�k"���SV?�YB��^[B���	�v��
i���ڦ��LȉP��\��r����m�C `�!������o��f@��EI�CA>84����<���x"M�`�	0��z[/q8s�x9�e�ܢL�g	Z��̘n�:�C)��*� ?I�Qn3H��Zsw�C�LVTHh$ ����X'�S�s>7��&�a�Ʌ	�/�>�'�V��\ �h*U�e��w�׺R�m�@���v�x}�j�7�ˌ��b��*�l|��C��-��Pl}6��z`7nU��*zf�G����f���X�sa�-�\8�.o{ ��=�V� K��ε'�.��K�4�Ϥ\r����c�S|�����O#�=`/�L塚�~z��ЖWB����N�����,�s0�?�^�g���v�i���g�����pO���ÿ��u�6�`'��t��GB���ޞ���z�>׼�]�*�^z�~��1������aCJ�z�D�}x����VM�����!h�"L<vC`�/�w����O�x�q>b|?o�Þa�A#���5q���0(ꯣ�@GJ l�;`��K�H�"��A��	OzuA+\�T��jh�R)���Pp�YAM��{j#QNm�m[�ߊX��n�Ԡ5�]�]ZҀv���u���悠�cZ�6��&�[�u�^�M]*�E� �2����[��*�^����T=����?�Ы�ֺ����Y�t4�y���'$��A+�I�`�.�[���PJ���7��|����08J�p��;�:]�vt8Wn분�ʭ�Rʦv�Vl���CL�Y�V��L*��Z�#$+�h��nf Q��nL���T&SHA-k��C3���N\x�3"����0@��UդC }��t���\�0�]�3κ5a+����>��3Oa5힍QJ-��'_r��$�kcd��Ǖx6�b�,T��f�(���܇�*.
]��'��׷�-U���Ց�Q˸��g�R����=�-�0�$+�ċ��=^�u'u��\<�/�.���c�����{��{�� �a������ó�=���b��~h�?Ӯ�M\��0{�N�Wԃ���3фv�@��h2��z�,��#j �Ӟ�~m:����l��}p�q��_��K��NЏ��4+�E�]���Wg����+��~��?���W��e6��zj�4LמBY۱¾�]�>g<Au���-������8Հ6����uk4��N�B	��b,cl�(����
ca���T4���D�÷�V� �E�U9�p�7��N3��#]�7I��2�C��T��ʚ��z�?&K���\�Z���o>�
]K����w�U�F�^Pj�a��Jl��̫�3�������Ŋ!e�������~ר��_Vi�bk�|]�B����:Uճ�j+��/�� Y <���c�X:uv�������AC�$��;��=e�z�(�J͗xI1E.�-��'�ґ��wU���nʭ�+�G�x�Qn�]��
2nP��B&�	5�-�2�\��)l�n2����z�tT=��S��8�̀�J�T�p6º-z.�������՟�5��yEj��nQ`~���>�P�k��Tc���4�BgQ�mVhC��#JR�E�e_��e�Z�������9VlY�E���~[L�"����*1��O�v�J����HM�<�6�[呏�S!=���TOXDGl�ހ���׏}�5���I�Z'�nu �;a2.P�=CH?����J�@�>�k�?bT�N��o��	az�[�X��aR��'�9d��_6�r}Ԙ=Q{?�5�4�l���4�Tn�^3VƩ鴃��[5��x48hץ�ل��c�=�Ge��v6wXz�w�U����½��~R��HU�� �#�](�S�n��J7왿��C�@���Ɵ��IP��$lo�F�Ò����u���$.�1+a�r�jG����1���[�"����}<�8Ў�^ 2#��oD�x���t�-�i�l5	/5=Ơ��Ϙ�8��P:���4mnk��7�B���ζ�@��=��͠��6�Tjm�
mUf[���'����'��8�+�8�Ӳo� �Z!r�|���J��'�ZGp�$:}��R/:
)�@[���#q���kTZz��%�%"�EZD���9�/hI��B)-�= �rK�����:�4�sɌ�����p9u|��9u��?}�����_v�9�"Y��IeI�D�i����)$![	�Jlg�r3��46���Fy��i���X������ه��P�B�&�����CE�m����S�n8����*����A�k��Tm���b�&&B���35+��{\�Ű� 
]
��B�>��D��;�t�}0���Zii�=2|�����C��X����oxh��hH�����jzɇe^	V�|P�U`f�j�ޗ$�Bq���bS=:Vh��`�Z٣��*�\����aS�ʒ;&�>:J�|6Vp@�������:���3Pdh�>�=� �C�{8�B�"ö�Dc�F��M��Q��~4�Ǔv}V�A��z���Q?e�s�ȿC�Bu���Ll�)�;��w�wC���ʇ!�D�F+3]�'�`�3�@����:�i�~��nx6��e���e&����6�����JP����=�qk�c�~\_�0%d%Id��ķ�v:������t;aq���'C�� 5���t�ފ����a�o7��_%�߶��`�~�hi�m[ӭ��ZY'�SQ(ؿHz[Y0��韠�~^}>e1������S�Nv������a�=_9���Ox�eZ����+�_���q<�c��i�"|�O���]��R#Wǿ:N��)5'�����+a#�D
2*ci�9>��-����(e�{��&Ҭ��E��H�%�^ӎ��m��q��d��J#A�*Ó��>ڲ���?
���<Gy8]�!$!��;�λ���K��?"ZCВ��K$�Ű�#(M��0iCY����jY[^�n��x�4:~H|�j�Xp��nc%Vvd8<:�^Ja{{]��%�a+��^N?\�޸R>��Z��΍\�%(����R����%J��������a�3&�0mf���b�(#D@�M	���(�`a6��j��e���:�Y�^��p��_[��v�km��Q�F찵�&�??c�Oķl�R8���)����/��f���&w�ܮ�y�����Z�l>���څy>�(��ʳ��9� %@ڿ+�zU���T�[9Ke��Ʉ뀕4d���B�|Țb����ʁ�Y&pv\0�;�/�q7lz�$�'x/�
v`(�]�k��!���d�#��ǋ��C}N$)ص�;�yn��S�������dzܓ�.�w�%���!*@<g8x �����īP�z�X�wEHw�u���g�ϾfI��>0n��,�f�\T�0T � �w��_ZI�(.�)�Ы� !qu���"	�*�ޛ����9f���q�zҎ︙;�nn��_R����9�8����օ�!�4͊|�О%�P��T:��P�I�m_�M6�
0����!y�=m���Ϗ���y��s��;7���f���(g�ޑ���*�qk��,�jW��b�n4?w��iq�}�M��~�o|��o|���|�+��h���,"�/����P�G�C��IҾ.:w��8Ҕ�I�|��)}Y96�
y�6�\�Ԅ<(R�ƿ��/�A��!]����l��~���: (a��D����w��rǔ�S���j�A���uy�J��6���R=i����k̔`�֜��q(/�����'�#93��p�}C:�?6�fR�M3mĖ�:�fy>r�7Z�{k6�o^i���Vo�$�wn������i�ԐFA�e�
Λ^��3���8��{����z,�"r��f�V��f��c3z�4�a!��;FAj���:��E�π��0���zL2|WYd���y�˾�8Vā���,��e�[�/�1�h�y��2�9�Zy�$Ŧ����K7e�H;/����I��y����t�����<�m6�����6�&L�f�_�f؏4�_By�;���Gr��3EnG�|���?Y:�T�AT� Ǽ���\���pJ�8a[��]��<���\��y��Kw����@~�9���N�Ǎ-}�$b��_�a��1�cI(��
A�O���+>��,���X��Uv�I��3�!q֙�B��6��|Ϫ�Z��:��|�Zp*TzB�ϧ�5�킴i�x��|w�4���x[���P�W<�h��x{�up��raK����3�,�x�\V�O�:���HF>k�E�||������~�[�z��'��������?���_�����g���6s,F>S���ʎ�|p����X[G�R:�8o��vڼ��T��R6��w�J��~�$�t!t�[wc;ʖ�|�B�����y���آ�U���Ɩ=:�UJo,y��>.=Z�_I[���n�d��D�K�f��m�Q��-�Kd)�~��YĢ8zs�G>�Y�)*�6ߵe�+��b�)a�6�ln!�0�E>���d�d��6mn���%�J�fڭ���	��(cB������x�����~��}mp��es�	� jcC�r�Fa4�$��S�v�� :�#OgQ	�N1Jߝ��.P:ؚ�(d"�S�?l$֫NlJ���_վ�1u��F��
����c~�sH��(�Q�[��+nh�eBD�1��&3��3@�<���'���[6���%����!fs\��9"�3�yZof��/��о��Or�;'u��۵�a��YH�HE'c���#�6�,��#�+�t�t��2{}��x�"���sG=�Ҏv��d�Sy��������t霧[ܰG���à#/���T:~]��1q���k���a[k*N�9���7�J���̚��h�B��^U,����N��C��]�������o��k�D�~���oa����C��-.�]�meopK����Xyk��;�ɟ�@�����/�R���3�>��W�������=ml���w~G������������������ui0���{�Bg;~��%��1_L�YM��;c1��T�2�!�m!M�su���vp�u���k�l��ȧϡR1�`����P�؆���a������d?a]���fV��[?��$b�#�ɞD�n���*l@�wd�^͊7�9@s�r������Ep?i����D)]�Gd��Տt�yݿ������e[��N��$���|G���Qfs[wn�����5�{s�����S=�����b�|�б���Gg%`�К!;˭CS��Ccp=�tL�+�;��DnW���;���h�&�N"n	E��+�I��6h)*T�8�<�;�#�J��?�]ɧ"�g�X���i�sN���7_|�x��ǫ�/�}h��&�Km^�<������?`���y�qI���?e�g��C�<O�we���&3/勓��=��8>��y��(�"�����b2��i���6�>RɿZ�� ̅��9�Zq�+}{h:��I:���fE���E�/6�fő�/8�v��z/�%3|�X˕_��i�<)BWcGrĵ�"sKO���d����:�W�:������QZ�>{Xl�a�TS������ix���3ƣ,��|����_��6��2}��x��o����	a�}��gsu��0��� �!]N>�Rh����B��5�/��sC=��;�[��/�+冚�O/���w}��-|{��HU�\����H��';ܩ�1��I�%i��4��F��#�>B2wUy�Z)blr�TC/d��'�~��{8W�m�aZ�(��s\�x:o`�OL+�k�!��픉��<Y�Ĳ#�$?(���ݼg��A�cҞ�Y282�i�!�8'�H���<�N�Eǯ��fHEV�f��k`�M��#�N���D�,��6!'��͆�D<���S�\$`�~�����|��F�]Oh��Ͷ��Cܕ��P�-�Rmv�׆����1mpuB��7�|	����7����g_h�����!�7����mh��&X����7��gL���[/�۱$�=�۝�e7$S2�8�����U*��cҋq�q�>t�9��л��_��ù���)��=�z6��q.�p��9׃�Y�Nrk|�yG�L�.�}*�D�38�M�M�+��э�wn�\�7ȃ�9_��0�}7Lu�y�����P
����^i��*s�;�"Ǳ�Vކ�p���}V����=����<��w�f;�M�������Z�"S�Q��wx����ˌyn:���&���?�u���]#>�wp}GO)v|n[��q�ݏ�O�TY�s��Z���b��������
����ò!=Q��{r�H���n%PI|+�X����D��q-��⏺]�{)	d�f�6����d��i���CE�x?�x���Y��1�:bh3C�q����Jt���b�W�e�I��2>]���Y�8{C��)��[�j����0Y����������ߤ��� L^�Nu�ᆱ�k�$;�uI�;�l<�#�Y����9��q ��@�"��&WQ�I޿N��e���Q����3���)�lŕwh����ŉ�jtY���D� (/㎣���wQ����'ޘl�ɛo�9�����C�6�(�'�z!�y��Lw��{��i�6��T�$�4�ښ���AW#̋R.�!��7��n%˵��L�4���/�!����z�HH��g�G�,7�3����%c�v&�K÷�J�1H.��a"֫<��.=���Ң摶;OP�M���ʴ�����a��$���
h,���^{H��e}n���q�pp���|�Ad�����)�$<�R�!��J`R7t5q���U��G�8���)���g�t����������N�7���+�~�t���ebo�G�
�m�d��U�G�EX}a�gl���������������s�����04)�TL�n�E~A战j4�������G@���s���)����V���7y.���:OIM����H�o�x�@������c����F��0�d�+?B���7Ѩ�C3i�֛��z3G9kPw���[��T��$s�o����P�(3nH<�8�_)��C�<������[o��i���ʘ;�zF���>&F���P�?��> {#��˫��g3�Y�>˱�g~ɾ���ʿA����~��~��{�y������}���ڜ��yæ���vv����kyզ��������R:�N}-g햪��17P�,��D�-�6}�n*��`��NS���=6���|.��Ӊ4�	�4y�<!*~:J	�/Nt�y�� <��W�9&_��A�#&9��d�wp�&�m��40��M<Q�@ރ�r�F��!��[�ԅ�4�LB�N���������Mji�b4lO'�/�����:.78��`!|ж� ��J��>!RJu�ӱ��b���}�`���/~.h~�{c�+k��p�^p���R����.v%�d(�7��Ҷ�����gޝ��K}�Vyx����l���Q�FWb�z��⎭6v�ʖ
�9t)sKI�=��q�pJ8Wun�qc?k�K�A�ֱ(u�
�F\��5B�Y������h[���j[��sU�C����3��x��K;b��v�g����k?�o�)�� �r�葧��Z�d��v ���
o/�G߀�����h:i��	���)eNb����������o?���o?~�k_{|�ɧ����������}��g _��S}��8F�!�;���At�[�Nu��*C�v�F��A}�jgj�JֱO����,Fc�r�9�]]�>�o�����V���2>�:Ȯ�@ܜS
/7�x4D2�ᵦ�X�;ol�U�I��p��U;����ͦ�%[���u���3^c؟�#	ds�����U<�����&lE����ݟ��/e�󎍫6�b�{����WxFv_��7�W<6��g��>@꫗*Gk.j�'b��岬��w˪�_~L������������~��'��}����?x����_����j��i�F'�C��l����VNxW����P��B����kr3��w"�㍧:�͒��c5�ߡ����_�eP�]'��A��������srx����ń�����G6�lj�S�=1Y0��1��P��I T"ʦ�9t��
�?����0�lA|<�}���('���'��F����k��5/��Ft��m�^S�:�vVJ��!���@ݦ�X��s�	�_ھ�9y�BjǾ;��y��>|Nh^�]��7L����m�F�jC�B����aa�8���!G�D<��!�^�s��o5�<P�W����^Aݤ�M�z59�f��׫��Uc������O�"B�!�X�j��wr�Kf�s�ЋYH�X8U�˛����0x ��;$�Ν�I٬FEw�Ԫ���x�݀��2��'Ŏ����w{9/���%��g�`D�)eFe�lt�yY̾R��u}���&b�v`�O&�`��Dʌsl��%�l�pBZݲ��k�@y_��c#��*7��y�<�^}��I6.�c������JD�K}�[3&�U��9�X�KGFbw�Z7��7D�H�A��MD߲����2M��2ł��Z�p{�hN4�+�)oȨS���sI��JZ�죄�z��w+��j����>�M~��} {���3��&YB�:eӑ2�س��#�r�C.��m|;B��Y�8��՞�6�޻�:�]amX���T>��٤zo:_�&o�^�߹��~��7�E׸����^Cln�O5s�>P_�T[��~�ײ�����㏾���W��ǯ��g�_���/���on�E":Yi�5c��bC��8v���t�|f��T��ɢ:�%����Wb�D~gBw�{h���ͦ�m�������G��#� �P�ޏOp�jP�Og�0��3�m�>AZ�ؼ��ړ�J�m6ڢawz�M� 5Z�	P��p��u�OH{�p��B��Gl
{"s��#�!i�K���z ٥؈s�s�VИ2ыߙ�~���-r�EG�\u�t8���7Z�1��(�P�t���9�Y�B�@��#�M��ſ�e�������	x.�}��y���%"m�r�"��~��o���sv���H�]�~�Q�zj�O�R?�&�MuQCO��E��d݂4�b)���?yO
�1:�=��ڢ��:'V6h*q�8�t�b&݀6{M�˱iǄ!��Z��sp�tps��R���_*���3�MER�%�+��stb���q?��D��Y�e'��<%�r�ao�-�i&��$�Ȑ�:��F�4�B�@�; 6�K1-����"�o���~�$ }mB���"G�ռF�%�Y��R�Ĳ�p?�ʻ{GΑ@�')�U �c����K��o�v[Wpv�*��p��q�O|��sE��9,��pH�7��K�1�>�����i�/�գ��(Yt�_i��:	���2K\⻧��:�-�=��	'�h��wk?g�'"w�1�؟��m�y��IF��/���"�[����eG����g��}��z|�����{���)o�e�>�H��ecs���Wڦ}���6�������{�_��O����js�\�sS�=�?&�6����4�����ͭכ[����
!�N������?m�wy��]��?һK_��8���ʦ4X�d3��ģc/(r�M�7�lrk!׀��z�k}�𛉠�����ز������}rȢI�}�v�T��'Щn��Q_��'�Npl5�EJc��Q�D~����y�u?_��y:Ɠ\�C'.+�X����c-Fc؅Ծ��[�B��e�/ܶ�	Ǭ^���T[tn��7�Qu<�4�N�mlP�2[�|�T�b'�2^�ƪa9t��q�x\�%��Ա�һ�V�6І~�п��1�u���T�Gy��/,����c�Ÿ��3N�^d��֌�BYy����C�E��-Z[y����H�Juө��`p�P�>��S!nÓ\��ar������Gƣ�6�_��aߋ�v��6���ݞ�tYٖ���G�e����\ԑ�>�xR�?�,�k��]eo:_%[��2K��d%�|>�mY�vj�n`����}$ʉ�����j+T}[���Q�b�+ß-���T���\�G����י_��z���U�n��8��K�ҡ+�A�8�������!?�y��}9H���S���,��C�V h�>���6v��?7�GK�{���7��e�/<���Gu�v��M��O�a�38��X����g⿡eߗs�:��s�=�(�i�񫍭����_����/�lp������>�����0��}��Gcs����{R���\q襥[�CT)���m=����O{s�7_zB��	m'9�cT�Mm��e����F��˼������1YSpY��`���Umn���]�K.�d�.��m_�;�4�6�SY���V����>;�[6��-"Y�>�(���Dw�Ik�("�s��J���U��6���a7�����t�O�]]�H쿊'�u�$���z�5W���w���j/Sܮ�P��޲�V$�}�i�3a�4�t,�^D�����*��Q/ڴ_�R��}�����-�y����0.��n��d2��Jy��M!2ø�0����b���'�;,�s�ֹM,zqa��I �z�F}�M�]��&����y�ج�a��C���&~��7�"�5>���\7��w�aC> ΅�W��R\��pZ)9��>*s,TG۪�t`�73[Xw�<��c��	k�؃�3y,O�>p�1x�_��q�g2C��e��6:N�����~T���k���*�$�1��M7�`+�۰~�,��X�v]�N�?�)r���iO1$+��"ʦ�=�G���'�V�=
��k:�㞟��kL����f�[���-��KU�:�ɹ�������=��W>�vO��\���*�Y�G�+N|���o���:��h׾Nhm�'͐��*���� ���g���I�>d�>��)�ڀ�a�7|Hx�?v�*��~�g��R6��}��-OB�D���V��~��񣣴O1���as�}�nsKF��]n����_js�x%�+߹��_�H�fs��us�M��3ln��#�c|^�[6~o��R"X��6�\@^�>wX��s��L-����2�tf��`������:�, �����߃��(��ͭ7�D����c�\_��V66Xvt��6<�݀N'\�>����� ۴}�:U ��R䝹 ��/�XG�]���l!�*�1��@�'���
��O!��{\T�	;.^�a��3�&\d���3��B��;��RA�F��}�ٙ ��F�ES9���l��o��ܙ�0R�=ɯ�|�Ak�Լ����8���Ms���8�sb)doRj=�F�7�ll!��jcÛZ�7ᥬ?�/1�g�]fs�5�/��1gMγn����4>{��l�>ep؈sڿ�+�%!F���ܱR�k���ɑ�m��*�	��z��Q��8����� e�d���`���e�O_�J k6���w���-�JQٙ�O��%= _���i�m'�����ʩ�n/b[c$[��s��؅k�:>�<�934j��� I;<�vl�ه�,1lUv-W�\�1Ub�U�����,�@�:2� �3��(~LH{,�p��U�-��`�b�G2ae�|Nk��Oٳ�Wݖy�:H߄���E�"�w��a���-w�y.ֿL����֚�������J�Rol���������j���-{7��_�&�[�dt�������p��*6�܄�>!�l�YN	�x?�s�O6��˟��[6�/������D��m���>�ɂ�@�B �D�Ə%�u>7��_�Vǻ΍�d�q�lD� bN �g��3�I}�w;v䮁�7��IE�I��Wcq$�����9=Q�"�R׍~^	�=�-~�OUl/�-��B�\Wt8�G~!#��G�z�_M�OW���D�\�����zOBm��P>��8��96-n�]�[fOh��I�>י�s:���C�,[��Z��wL��:���U�Y��}q%��;�W�@��z��vi��B�E{�E^����y��/θ8�L��5��&v�D~�L��C���j*?:/�z!%��T��k�o� ~�xs�Q���_��K���R�L,P>}P�Sɏ���NZ<	&k��⌝�q kH��l�ɤ��[���Eq_���#��U� ����[�*/-�V1Bݞ�Ob����G�ߡ��~���7�oDՇ��Q1�D���M\>_]���S�P��}S��t0��ڴ��b��j뼶�\v�����j�������١b���պ��A�<�й!�~(��7~��7�Lȡ�8���7�}���/&��d����|��k"{?��7w��j�%^ָ��ᕻ�b�y~-�/1��|�������lbeK1�g�K>s�<�?����B}��@�s`�_��O��޷��η���o7��*A�ڼk��|lp����-� ��!�\1����b�<���1��8d��R��YW�1�\��;�WR�t��{�h͗�������\�]G)����Lo��y'���'i�l������ؐ�On��y��i�'`��U6��{G�X�a�7X�Y��u��۝SO��^hŵ>��s5m�*���M�z9�k�����9}N:DӉ����ы�\�yR֔^�T+��a|��M��c��Gd��{�{/��Moz�M��]�͋��Ɩ���,`m�|QY��E�1��jg�){�_��b�~��T�F٦t��[���gU�ؐcu� =ӌ-��g���G�P���kQ}�X�3��Z/��k}m1�k���H��:N�J�ª��m�	�C�mCl���(��u8Q_��r�^A�i�_��L��y��ڼ#�ZoWg#�P]\;��8w�Q.r�l����8�T��F(��H=��I[�6g�W�W_N�:dA��Q�Oec��~զ�w'�E��W�	ٶA�^'���,{��?&��kN��m7�`y-�,����<�nm�RB�"|�ڟ�k#�u-�aٯ������U�v_�3�l���a9�kȹYk��v�#$�K��[mn�����c_�*��o���[��M�m�G�c»ȍ�<RC~]� ��e��.�*��<d�`ʇ�Vc�����ȇ3laJ���B�ƶ�.'&���6����2$Fe�?ˤ�Ǒ��"�M;�Wc��@X�N�z��(���#��#�P�z,�F�&/��u��փҍ����Y07���V�G(v��Zޓ�W�mk_ſϼ#I��N����/��~���Zd%#��QM��;2��P�k���JR��S���W�/Y��8�8Tiމ���z�����\�r��?����9�<�����/����������?��@��b�E ��m���5e��ѐ��C��v�36��*~�y���H*��Z6���W��.���#M�a��א�Y_�؍��%�XH�����qnеMȄ�3�m%�U� _"��\Ի�j���R�y��`���\���
�u\ј��P�so�TT�d|�����#�t<3i��I�(?���_|��b��A�s\k?��j�V�mh]���t��F�6�/�ve����{k�0LQ�ڎm�r���0��C����� �FO]�^Q��d�����*{��[�ݼ�D.�	��pl+�7�lcsɗ'MllY����@^���wkk]+_>��Wdy'Y�_J蛖l���[?ˋO�Ț�G��b�a˽��b�\�=���i@���*^?ʥ��o���6��u����G<:�Hl�S���6m!;��E�L`�B�!$xN,���2<%�V鏋Ϣ�	�S�v��@��������;�����b�	]�"0�?bɠ�Ej�����&l3��OY2;q�z�#������E�i�j�h�@�A��ms��E��+�C�19
����.��B����/�2�D�h�ټ<���75{�����?S�9-��5i-�>\q��Q��Jj��������w�}���ٙ^�C����r��̝�-OS+�ci������p� �՞�,ȴŧ��;\�F�7(��*"�-���6���7>��G���n�xK�^��o�w&1��4^%nvL�K%�o��2��ʧ�$Z����#�.�%ѱ_�9�ʂ�<�LfL;�JD;�5`�塍��6&�˗JCo6�1�-�>y.� ��z��|&�~�g��m]��g�����j����?�ה ����|^F�H���Eg���ʷ�0]��ȸ�4}O�sT�k�ؘW���*ق�+J^4aCI�;6��T�c�U���Ǎ���dH���E�����ٵ�Zq�<�Uz�B\��i�=�7Ԏ�?	x��>NX��7�=���w�;Ȭ���6��C��N-���zE��s��:o�%?2�wUǾC��b���Un.�O�őǌ����T7(����f)%���\�@��<��B�\K���~glnY�L�+���@>�Iٷ��	8�v<�5�4�H)UoxQ�Z��'a�*��Ρ��;f��"�[�E.�����+ȶ��^ f��c]���O"��ZH�-'n�	����j@�O�Su��Q�����~���4S~�]��� N�I��w��	�V}�r��DH�菼��|��j�7:���	�����Ug9�)d��̠��-)s �n�6 s��il���o;:8��!Lؓ���|���sZ�ŧ1��!A��C��V~�v�yag��eN���0�Q�;���m�yji-wz��y0R�������[,�س�J�a�s��D6L���ƶ��mƈ��G.�h�\tj]��3ƭ��)kll�Z*�EYe�W�ͼm�Gd^ˉ�:�K�*�/ܮ[ϻ��>�W�����5lYe��oD���°{���t(2+y#�]����۸�G�@�>9B}V��}%�8�����q�Ժ�I��o���}}��B���H��I��P��߄2�Qi�躅r�(o�3�*T��J϶���L�S�lj`꘨g�#��dol��d��}������&�B}��țZ(Y�3y��X��$�����S+�xG��KR�q�ͳ}���oLHs�����j��>O��o�_A�0���X�����V����U��#�v{���J�����k	|[M����aC&���/F5&4��:�%�����[&���x��|��]�@�+/e��E��,Ltz:����گ0.TG�o��G����ũ[��/�i��qE����ցo����J]A��ң�A�(c\(�'��I�~�H)�e-��2ᗰm���9�(V����r�H���x";��㱹�`����]J�ԟ�Uk�.f{�p����wz�*6H[>�j��cA�H�#oU�N��^�Sfl��y�"�z��Ӝ�GPF;��.8��Wz��?wp7�<s���/c�P�ݠs���r�v\X�ɼӹ��Ҷ�w>>��-oj��0GW�Yw�xM��2k_�0l�n�S�r~�&�l<���"l�OEo9�-��5����[l+v�p�k%wB6$j�R���^֍"vs��t1eٌ�2Nl���J�<A��$�?���o�@;I���dU��F ���!�|�i��-�^�g�(�}��2$,�[��C�I�φ��w�0q����H2t1�#��9�(��Ƕ�q>��F��u�XFǺ��#�o�ξǸ/�E�DiǸ7u>�����9�~D�[Ma�q*�s]��H�{�����R��Ʌ1���/ko�:��W>U��uqFh�%p���Ῠ~]б����ϛZ�~�Q��������@{�%{En�z��^c��6�S��y�x)���P���s��~�k�X�O>}|,"����������-�2I�L�܌���䱲�H�s���?��7���?~��?{��~o�BY:���MT.�G���|S)0B�b�2]S8�tM��6���D�-�N��97R��w;�<�eڃLd��2�3�����h�:����o﵍�}�`�?mH��U�]�W�Lo�m�>,{E._�H-g��%�ɒ�9�e�t��������O^����>����f�Tvl'���WD���l�L�e�_��h}�:=��Z�(5j��]�����R��m�(¢7=��T}
)W&�a�9ܞ��F�s�[����y�ͬl|L�?���ߑ��\��غ�9OX��뀬 ㅿ6���AZ^�WF
��ŀM4c WG���k�G����H�M���M=Sq����АT�s'�tY�΄�?c��=����^[���Qμܑ�,3�w�P�:Mծ���*?��c�w����S�T6�N?E�:�{�Qg��������}��}�\�;��&�Nz0+��2Kl ���5^e&~T�!=Q�V�%g�M�	����Z�t�.=C1���mWU��^���B��*4��"�dcP�P�\ >���b\E��Z�ǆ2��BZƲ��0��י��!������lR�;��<Qml;���#�>E�n:~�Z֦�w���RI؞��A�u��7�bcK�Z���žP]n*d|1��kņ��@�{3I�7u�Я���������B�&W-��X�ƻ1� �Q�S����X:��ˀ|�#-
lE5��p-�����V��k�v��ch��lp1{�.x�����VQy���P?���K�'*������q���)~HM~�����O����k��*�Qr�|%�⏺������N$�z��2'Z���/'�x�/s�E�	�O5|���_�iJ����f�OT�= 1���I'9n�z�{!Rj�~�����K]�r�w[-:d�Q<���]�C����1}�i�Zɾ��]�B��B�����EĖ^�A^$m���bld�o6�kߌ��佱չ��0"�qol����9�`�%��)3-[�!�m��#_�c�������	���X��/���O��M4x+[�\��,��3����h���Cض���Q���59�S�C��!����E�<�i����9�L=o|�!�t�m��G�;=�c�6�����w,�Nj��@�?�=+Ya�M���?:�vv|*�Ze��y�ˀ�`C	ɇ��LHJFu_�ƞEL��5����+^m��q�u�"���T6���C~!|���N�n���s���/l��ĝyG^�خ �[pZG��]7����b�P�^��l�|r�8��c���^�,O����iݹ��E5z��^;���ؗ_��w{U���;�~�9s�!���?$]�K�x�ľ���Pʗ�S������/���v����ʾ9K����H�;'.9�L�Z�	�����H	�Q,�~��gY5 ���a٢���Sdþ�?^4� �O��1�81c���Z��D��t�[���l���W��G�|��A��;=~�������a8^�P��|��q=�փ�tBۼ�}{��W�$m�K��1+i����l$g�O1yf�W���ڇL����l(K9� ��]^p*��0h�`�;��u���"���8�i��Tpb}�[��w�iH]1۱C��I~:V��^ԏ�qF��^��/t>i�c�Q� �.��q�䰇�<��8K�+Ҿ�OdDn{�k�	?x�Q����͹�s�� �k?��Gv��N�X�Yg�m. u��CS��5ڑ|���YwS���1w7y���g�:޴'bA���7!����*��u��92P��,�  �7IDATKmjy�R�]Ҏ3Y�69�ɷF���٠by+pR1u��?�c&��|ڌ;ʄ�B}�ێ��xY3E�f;�˹�o��l�EȂe��5JW����2WX����Sݡ�X��h{�W��(�мQ�����@�n�d��S�1w�SQ\���z����� ��2��w�ې�úƆ���"���s?���w+F�L���ٳ�6������yl?F��sc��sZ�Nh���~��8Ģ����,���%�(�8X��?�Kw��ԏ$�m�ظb,��NĖ��.��>�S�|C���n#O�&峹�LY���$|<I��O��y�7E��@(ul�qH������^~����~����8����?����V�!� gB�刁S����Q֢$������O�o@=q�	�� x@lVv�)5�b�md2��wT���iܙ-Gh�Ḑ*e�碀�ׯ�|�
���dbR��p���c�>�Y�8�>���]/=EQ�h���
�'M�(+~�z��^6��K�%�P�gp�³��[e�N |�����oI�O�K>�}�Wi�5����/ڇA��6YƯ=��\�A�h8��}in0��lk���%U���Xm����|@�c"�U>�Y��?Q�8f���|�i�*.�W�����T�P��wGn�oM֛s��~���Ҧ�]y���O?�][_6{,�,��}�C��ց�Zx֖7��)[?[��wl�`��`D�㼎	�.:�K�g\�4gM�9�Bo=��7���1�jv�h���lwE����C]���u� ���O�tne�/�5YI2����&����cs~@��u���xz|Y3����G�%ΐ�yRba~�~���b���cNZmX�"����l2��b�>֫�Z��Դ�/h�iw�ډ�y����X��j�t�
A2�C���3]��ϫ�߆գ8GyMQ�x~{���E �E,�;>S�oj�	��~�9h���q�:�]��"��U5'������]�y�� ��c�HY�{�>�u�o�*6��4zη�q��Q���/q #{�3>'�J�ӟ��lS��6!3I�g�p��,���I�W�Gi,��2lh��������K�_���|�#,M����bYa��U�1��?������/��w�������[mn��6�1��6-�(�Hf��$T��.k�F&s�]Hr7�#�����ڬ��650������$2@v|������?�-LF(c�%�&ع2��#nlʶ�h�3�6��>}�q��$V�'�v(�L�"�c��I����[��9�O ��CsuqSڶڞO��R׭�C��b�ٲGfM�8Wu]߹�Ķ���⩺k��*�+��ղ�H0.L W�����ڱ�t�B{���¾�7�Jq)�#f���X�Ë�,H�3�"�&ק�/��p�ѤZ��\߰u|,�G�:0�/��h�ј�X�}*a�5��)�ln��%wn�oz��Z�g�����@<ߵ�\�/�y�bè�%_�z�Z�Z&dÙ8��}թ��k�� fs�kM��~����E�߬����2Oߪ��7��?��J��o6��?�D���o�}�c���)q���|�yU6/��GD��<]ۆ'�v�W��A����k��n���P���u���c��wjf��O�jt�W�A����]g��8/5>?-@]��Y�ʟ��a6����HY�_�6�Ts�D�	u>���i��2@��*�:�����X�g���wS���m���������䮵�w�rZ�Ք*}��c�C>�sn��@�%>��)�L�;�;���  @߿O�>V`�-/��/�t�b�T����W�ź�v\��<�ћD�6��Ew����w���/��_�}���7�f�#߰S�𼾩p�o����D��yS�G�i�`(���=����1�ؼ�-��U�����O{s�smn���7_r�6�g6���#N\��;ˀ�Og�X�m�?u�7��A� ����Y���$7_(����/ �	?yo|yd�.�QDCi�����O���{�D��۔�.�V��]��aB28���۪W6�'>t
s�ݠEKd�g�J��F\~)�G.�;/�{�Y�:pl���Bz��⧗��/)�g�T�v��|R7�C?}A4w�T&{��I��+�E-�|��R3.��1�<�}zA��s*�XU�uU�1c�&�ȷ�D�]�gxQ����k:�~��]! �:��zWH�Ʀ�g |�O���xz�@Dp��iL�X�?|T��ݱ�A����p)3��I��_}��e�*~8��؋��SF�_$�f�Pk�m���7���z�Ϝ��#V�YQr��Y�EρN����X��L�]b�'Q��7SH=��I0���V��2���p�Ô!Vg�Hv�>�a�$|]w�w5���e�MSn�痘��8�5���w$��r����J�n�,�O���m6���Q�eh&�\�t(��d�p��x�1�ґ?!���E�Ô�:>�.)���eo�ʷ�� �?�Q���8������z�l*���#?@M�E��j�`����[T㡑Q
q�1��gy-�j�?����*���S�����S뻵��eo�x��<���7���������%eo�R�1GX�z���ai7�9\�\�'n�������;��*z��P��빠�0!m~I_���	ml!��~�����~���?�ß>~���}������|��֋6���Aˠ�e˓��r�/u� s���Np}es�[��x��OY�.�b�W�{"�#Y����Q�u�?���r�,},��|��o}b?�� �"g�M�Á��Li//هb�ɰ^x���v�m�_g��e�P%m�\��'bp�\g�]���'=%���_�w�7�r�ؚ�q�8��San*�˽XSP����,��dɠ��ڤ�/�)J���PE��;�ԭ�4�0��	�
��{�Zm�s?�xqt|��*l��������o�ȓF�>s���R�<�;�3� ��/^w�D�W|>1��v�S�\�z����*���4_�ô��q^+��|�7�ܹ��6k~�綌����خ���@ԟ|y��Z��T�)��b�p��▸�a��U�d:���E�k~+b�m�Q�.��\�1APU�We�J�/m՟��tc�(T�(���� ܎��:�z_W�b=�x�ڐM��z�[�>�4�����R��|R�1�n���t0Ŧ�������N<0O|�&����No����7���s�Mh���8Y��&7����~qȇ_T�����<�m���ȅU�`�.��y�`lElj?��\mnً1k9�R��߸d��_�xs���[6����H����S��[,c�����ۗ��į�'N���Z��X��[��o�����ؒ:�ZOs�@���r1��i>u#����}�e�3i��~�P���˟?��~�����vne��IV'���'u ������� ����͝[�+@2������� ���!�`?�w$,˺ģ	�A�G{<A8a�+Ŗ�ǅb�?|�W��j3��ɘ����0E��w����(�J*��`L�dN�"1���,U���U�<�S���oW �h����w���z���%��y��؉��T=���T�����N탴3?s�l�3�rb'TN͔=�T��-�F�?G?T989Q�Џ�C�J��"[i�O�J�!������<�F�M�߂0�%�|N�ys�9������;X��8×�1۾��9�a��G�x��GݬYZ���;�o
Ы�&mS�:�y�E������~S_k[bF<}r	{��o`�r>��|�	�}��TӋFjuR��	$җ���f�sj���"�C-n\^�*����}���`vm�ܹ�|���g+sQ���b���t�<����k3v�7u�aM�u���`�%�7e%֢8E&�$��"��6����p�,Z�`U�=h��f.��y��T��80S��Fl�#��N,��3��/RN;�� V��<����k�������J��ν�:�]�R�aS�:�i��/�\��S6���e�	S�?��0��w���_7 �����gh�h�k�q��0�mЁ?�;�7ה����es+i3�9�bc˗�D/^?^�~�o���/~�����m{�,�.�N�����H@C�J�5
��G^ҙ�)Wn�s
&yx�N�4��O/.\�E�����}�]r�`D���&�/��`1��!x@W":�.����,�K��O;g��+�U��^4�S��$�_��}�&}�Du<��3k�W�"�WQ�����n����dR�}@��)*ȯ~
]�U�	��6��]P�ep6P�O�3��:mkǾhSW�e�� i�>p��r$��k��Te��j��pMK���ل⭲�{��Uq�"^�[�.H��3b�s��;���|Ta Ǣ��<ֺ�u����0�	�d,��S9�fr���&qN�._�����K�5�Z,I�app&��WU8�Ԁ�	F�Fڇ���|������5b&�bڶ�%2l�M߅�]Y�@U�fx+<>���b���^����[���l�!N�$�v���p�t�6��6�6c�ͭ��+�8\��6X�-�t��D�i��n�<we�U�(:.�+\Ն��������� jU���>`E\��u��3�M��L�*�V�)�� �u2��� 6�گ8�x�ZRD�z��Ǧy���#{ml�8|�f���[��D�K�d֝�H[Aƃ�����<�onUiiԥ��U?`�9ܩy)�94y�ϋyRr�v��o~R�<s����Ý��c	"o�݋M�H繄�,�,��3�3�R�u�|*�*�3?Vg�݂�n$��^P�:#�O�8�͑V]6�>���������S���)�ǅ��:C�i>i��c}rP�?��g�HD[^8��2"cd�`?O���6Ά���
s>��: ����V;�ŷǫ��I?0<��;;ɹ?�/���:�V� �*~�CX˝�nң�,�U�X�v]s �xU��Z�Ե�Zk���z[�1�FO�~�3���]��^lK�o��q���a����}b�T���j�����
�瓋b�������vVۏCcni|���lp}�6 �/;�z0P���Qp�T�u�7�|Dȯ2�&wn}�p���R��x���1Pz��j����:���Q,Y�tG��1V"nS����r�ر���'u3/�嶷�~O�7��k�|�Q�l�}ڈ���|�~c�,��?s.p�{�-7O��=�16�B�{��|+����N�&��%tnǝ�����}�;���?l�Y���kݓ7lo7���i�2�cl�M9��:�rB�5��XD:�}����?��}X.DB�?���\_���Zã5�/͓Z���7���f��9١L�ыXY��g�摄��r���s���>/�}C���^���l��>d�	��RrĄ�^�㱙�������js�������?�斟���VA��q^ྫྷ������M��.�G��"�#��eD#�x���BB���PS7ʦЏ(>���<��^e���Ε���&ͷ��t&�4m�9�A)m! ^tiþ�J�����h�t:��a:{��-�c��;�2��hٔs��l��:a�KVe|�!O��&����ǝ��� ��	:�s
��\���G hᣁ���/���Nf������R1j�^a�������Z`fҟg~;������Dc�v$�/�<����{�֏5�n�`���ǴM|�('.�zY�d�1k^[}^��kه����?:ǳ��7�\ X3d�;!^�*teؿ�B���y���:ܱ�O��9J���I�Ưo0��~����|�9QuƗv�n�-���Dn9�V�8R^���1��=�\���Z��́4��f)�Ŷe��D�^� &c?.�a�� \� ������ʭ��G&c���G�\K��W����gf����tc|�n�3�9�t�|�����7"�h�y�UlSf�CeuL1���?��7ҿ��jP�|�/�c�6���y�U�#��� ���|�?�I��l&!��8�.�oYR�Ĺ��WcΚ��D�kT�OB)����|�y��\�7��z�ŁHNy���fis�TsQ��D�{=�O��/�m��Wr]f����@��NPN2�ZO��ծZ���~��6�}��g�s{��b&��!��
m9�/��w�k���|j�;W2��a�����	f�����N�I2y=ٜ�~��>u� t���z��v�Tw2�ܖ��P_��V3��dVm�/�.�M��
Z@�?|4s�3�������IQ��4����
��a�6��
�JĢ�|�e�>Qi��zs+�Z��̅�q�B��R���@�C����#>�ZK���y�=2�>ZqX";�X Ch����@h�k4?ң�t��i`C��w�ӟE��+����y^�otP�X�g7w�3]�Ĕ�c�@jb����L�:�W�,U~G��"��A�S���X��E֋��,/���v|s^�b���_"Ӻ�?���kc��3�����!��Fr��uQ�[��.�E�}����#Q����W+`�%�)�-ִ��/�荤�9�k-V�(b_�E��gN����uߊ�;��	4�*�ذ&�ɻ�c��A������43�Y��E���A����ɩt������R�AáF�oX�}qp|D�q���mG��Q&�M��1Ō��y.��9綥�v�5�S,�
�����V4������T���$?Ǜqix�YkL��@dMl'^�՞�[�7�k̅jk݌�K\\Լ/R���V>u����&���
��O�*O�eR�*���x�/��k��a��K{6�/��jc����o���Umn����o��d6t0�Ms�:(�,'j��� (*�o��mu>�zŔ);u:�u�Q�����(N)
ͳ����{���<��C��6�T�8��;��e���f��u1���
�^�9'��I��XX��¨�U1�����29=BtW��(��}vҷzl$jq�m����y.d��N�S&�Ov��R���sֆwA�9	�bb�e��1l��6�I5�O6�aGX���=����Я�h�be��uH�c~� KE�����J^dYɶ�s�A̖�ֽ(�VL�w��,�ܿ�$t��c��\�ٮH�9l�Cη���:�e#d��H˶R-ÿ����EF碿��>�<��H6�"4��ln�X��q(�Ɔ���S|�c����TF�ן�^�r���M^�SZ�tט���J�t^�u<��l�(՚�������\@��u���$�;�<t�I�a�U�1w�7ڷ��Z���_oh]=��y���@5Gm�к�f���-F��T�at�X��6��q�o'JΒ��]Y��o����~��������f~�4�O�зqJj��C�2/h����$��#x"�h�H��,��-5��-~$����]n��J��͢lK�=�I�����ڊ���N�����w!~���>Y�ʷ��O[<W�GʾN�t�u�ć�Y�?]W<d>fs+����`d�'o���q�@�M-��bs�gln��?��6�����_�7��;G���XC��+耬t�'���nP�lJJ&kA�N�?�Kg ������J��`9:����le�����F�2|iڎ\��g0�X�O�0QH�:�f#��pu�D�(!X�����j�t��J魨�9},��\�.��8:&'njb�]Nj���xdB[�}h�ȹ0Ѷ'Y����79�q����+F�K�/X�o�]%�"�mYE<�-�@ˠ{�<����E���U�>ť���V�:��yS�ó�c���V�q���h�Zp��M�Yy�������hs���'�M2�� \i�u{����>6Xl%�����|����=��<�2�6����,Q~z'�<Ȏ(�<o���r�#�x}c�ځxk�;��i[�hb@6��巇�-�^A���#����g�?���-��j��+��;�]lQ�tupK7�P��"��m@�7/�a��^?rS�2w'f�$B:�%R��tPWa)[�P�E�`��h�\:���b�~�d�#�sʊU���qmо�:)�OF>_�}-���k�yVՎ��6����,O�QvU�!�12��T>8TM���S�7�qL��ƼQ��ME@�"�'��4{H��xno�_�W�X��*�������A�5��HoPx|�L�Z�G��^x��+���mn�p�f�ß�d�k����~�#�����^����������������7�Pp�Yj6@+��Hl�;j���ɲb��~}��%ش�z= .�H�3´��>������0'��`U&��j�6�u�R�P�)J<��JV�A�+}��21��6[2F��݇L�ҵ�� ��.��Kw�U�s��?Q��I1v�;��٧]���<��(ְ'\�Tյ�M��w�<�Q�N6>ϸ�_a��䐯lڷ1�����e�֊�����Ĵg���}D�������$�m�å\$�P���uvSF�8?*;�`ڱ����Ed���h 4�kCۿ-���Z�5��?��7ٺ���/q5�X*�&��P�~������E�.,MCȂ74�:[�,ޠ�"���0�+��qlk��+9�+������uE��
��#Y����#5rO{G��4��?P�i���ƔC:,~I:��Ɔ��Th|}}V�2Eݏ�Ay�Dޱ(~�RV]2l����-ɇ���e�����]頒�A��m{�'c]v�n�`�/^ј��p���E�ŇAZ�a�H,�u&o���f��m_�0�qb]�?��#��[[�_�l���:7 ~C�����[[nR.yǨ6z]7D��v`�S�v����Z��6��V����ڨڬ6ġ7�y|�_��w���o<������֓�-�`k��I0Y��$x�ll�C4]�CXt	ʩǆ8���T����,[�cp*��S$�RF�Ԧe��B��F���˞�JG}R�VkK��
UV~��9⇲95���	5f&lA�:
�'6�[���J�T=��8�+�F˹�{\��!����4���u�a����f7�d���"΄�dG��7X۾C�_��g����`��b���,/�sAI�3���;bȟ)�2���<�D����?�8ɏx������9�9��]6��;�<����z���V�;� �yz��聆��26�1�ǅ��ӕ@�P���W�T��kn�l�
������.w�m���,u���7�f��|����hX�5v�o^[ł%�_�[S�\G��_u�Iɟ_;��x��Y��N�ۿ$��J��_�ak�K�y��g��tzx2ڞX���
UU���2?��?��mH ����C(�U0��Q�6H���"|�e�I��B��'��50��t8���oI�"0�7wl_�g���5h��7е��5�?��ZS[�������@'�⓲�u��wS�ԲѬ�'v��y�Ǭ�z2�{.M̓.���X���b�L�S��ė�����z����y|�w����7�V�[$��(cn\��$��P9H6R8+[E�C�|��yЋ|.�"�&|���e��Y��k�+��JlB�h�pu�Ai�H-&yʰ��yI7�ь�y��/�ɬ������4�t��۰��ؾ�_�Ƴ��#_)s���X�ioq�#�+N��:G�D�"e�t���1D���W�l&^j����wj��Il���u��7:=ÍH��\e���0NN�ˏ(��&D��ܕb�} ��2�U'�-�+�ϗ�8չ>u+?TP����#���:p��gb�^����w|e��Df,s^q�-[�����yc�����Y��-P5:3�J�e����"��1�>�EˉM�03�A�Zm'�M�E�To�����<z;�ɆoTo�E��5u�U��p��p*��:�}����.�׺�H�Va6>P�.�ä*{.A�m���\ϛ������j�1��9�|�!�j��� |%�A���{����y�+J�����S-ֺ�GB~#����Б�3��B��,[(��M�ni�E������6��ll�F��ᳶyC�u`�gК����9d�o�5��e/�,�%P[���W?��w��η����x��������ͳ���H�,���UaĪ@m���E�DE�`�W��n��?+��j��'y<�:�.Dt>Ie[�����g�h��j�K���ϒɾ�e�������|�.�9����i�P�a�%��c��|s�N�BO���g��;�`N;6c4mQ]�p��A
���Ҡ���3�=�W�r�M�FBڶ̈�]m�,�����e�Y4�b)��M�<l�]��j�҆�OU�t�Y��ItPU/.�W�
Y���zY�zٱ��pd
Sæ�r%z��[�a��_�~��<A&cuo�v���HYc���t�o�a��:���a"�ܹ%����e�u_w8�<y]��׵�q�G �t�b�YO��Vư�\��ȝp�5�=�"�o����F��X��Yh؆��8_��g2I\M����}�]S)��[���9�a�����V�Ys��}0���Ku@���:Cb��'����i�p��� �EvT��x]>��9�8����땷�m3z�R�������֝�q������m����!Xi��:;�Ƣ��{0�3�'��KO�[����躪����WJ_����չ��@>R�q���@�7�)��D�qu)/��ٛesd�������.kL5�Z㋱싴��6fKѪ�U�K���71���$}���=�ńW���>{���~�����?���w���@�gI���0Yf�\�k��"DR�U&�«c�+�ސ��r�⥲ڶ-��c]&y`{�!�(zИ,�ǿ����{Sr�|��<N��m���r�h���;R���E�:���q9�#�>KP���<7�~�v>u!M�晟r~�@|��,�|�������R�2�(/�Oc�N�/҉}�)ގ}����*�J`EX�����3̯�{W��A�\8�%4e��o�;0�ⶒ�T�����(Z��_�ߤy�Sɱ�\W�V��r��<?Z�ߞ[ě,o�!6��nJ.�)K�O����eq�_1��R�cX^Ķ�{�D�V�[}2�'|Z�i6z�Rfm���ޕ�p�'opW�9��%dΤC�8���><#��ǁ�G�}��$׎~>���?��j��C���[�Sl犰�%���ϱ�w�9pGB��p�����R�vmx�"�Si$��Q �\;S�I��Au>ys��C�h](�'��&m�L�U�j�Bbw��8'Ч�)"6��d�2�Jh�1��x��[~q`}�V9�hT~�.С���_Q�s��9��R�)O���3'�yc_ >����ڜ�����k���U>#�/�y�V�����c	tB2��mp����r�A������J��L4�s�U�GP�?l��D�5����B鉐��Z��/�Dv����Ż�m���/O�k��R���^/�𕱬|�Ӥ�aW�uNd������QN��ŀ˦c}bd¥�I@�N����?R��c�%����O�X�lM�l@$����>W����H�o�b�)�p����]�ݝu�{G*B��E�WW㳕�m+9B0o��Pn��k~�wr7�h��T��p���U�D1�;��\�K�;�g�/���v�E�7��|�� k^��Y|����{ 5���&^��B�]���܇�pxɈ�m�e�
��G�&��;�F�"k}�}�T�b�F�"Sp:�� �'5_Q?]̚��3	ZIF_\H/l��5��^��g^m� ���/��א�x�K�M]�!�H]�0�|/�T������Ч���>��+���C�ys���N���tn��p�>��Jy���X��Q��|sp�����s�r���wE��~6�՛=6zYc����T��n}Ak�ǟ֗��f�LyUG,}	��s�ru���mQΛز.�U��f�1��a�П	t
*��6��<9%������N���3~��_������~,�k���ǋ��g���"��j��J<���t]�%$Bױa���m=CA�E&;s���2�̝�����x�B!��:2�q ������Y��wW|�e�⮣�����'C�e��R����W�H��QȀ��o_tV�GbW�7�6DN]��~�u�<��~�\���V"�F�H�֭����]O.�nI{<B�9����T��J�`;���[/�57	M���{O��7��m��b�eE�F�F�l��3N����#�>'�S�TE|�y�2��v�[����XR{�3�)�d�VDc"�Q��l�;���m��H|X�v��b�Y��s��+ʧm�9hs��d�_B�w2�}�O�<��u����[�Z�Ie�{k�U�׶긬o�<��'���01��&0#�����y�#���t�#�K������2�׃�h[��˫�����{��Ya�~��P����َ�y�oz���Ʊ\R�
3��d^�H9|��H-U�z�f�}�����䇊;R:2��q@��i��k����/�7:'�Ib�m�L\�YKz=�5�U���Nm�;��Ō�mۜ����l��R8;�`]����z7�u�N�/�֛羛I��K��;��Տ#xc����+��7�bz��>� ���8��0I�~�_6��Wl�+�L��qb��� a�B�NA��4�8k?貈8Y1-��^���'+_��Ho~�����O��=~�?}���z����?q@�Nj7e�8uX���@z��<����¡�:�uد�C:T��k��R�!��=����V�p6����S>�߲�A�}�T��8e�p!z���@���1���t����U������M#|'��+h{u�C_3�K;��U�:���\ƥbY�:4�b]�� �xN�������;��*uMNY(J�	[c�6'X
��EFL.�${-G��䦽�z�"o�2�W`�6ew�����	� ���nH��o7�����I���]h�Q}���4jSQ��&t� W�f�iK����m���ic��>j�)߲�⍖5vf�\1�'�*"d�[���#S<���m]p��e1f�טi.4�<Z���e����+-��#��5�/n�܍�{-� y��rq��>�O�o�y�w�
U8F��M�R7e��k��S��Òjo0�L��l4���
�rߊP"L�!��&�U��x����6߲��-v�:���Xj�
���ΐ�,��?S��'�`��v�7��Re��K�?]g%K�\E�u�������]�!�YO~L����863f}+��2�f��#�K1�~�T5{_��0=�6���Pw�z���l�M�7�b1��M4��Zj��V]�'T���cO&_ٛIO<����"~\i�Q��B𼓍����NN�<�*֊��	���)��f�������Ԇ�?��������������6���oi��!���ܘ`(�ܸ�����R�Hi]w���n$0��R�]�������H*�������9�e0�����փ��^?�Ə7��@�_O�D�~��Γ��D�K01
v{��qD���DY��c5p�X��p��Cw����*�N��;����R�q�'c�w�ew�b�<ʧ���R����l�s��[ƿ���֑�%��8y���8�9� gIM����1��[�JR&�I6�g�w���y�c���3�M<��:�f�WW��x�����Ll7�޷!�]�9*kp8"U�s�\Ѷ��&�O/��&V�a�7�E��-�z�)qt����lp}���^�ks�a7�\2���|D8˩z\�'��v�cuT�z<(�/�O",1�[�~�͟Q�{AM��1�c�oTQ�(���c՜���aD��6Ѭ���PY7��zYa��+��Xl'2����C�[��c�a��A�ٌm����!���C�u�)�<�-[1�Bi}�u���*O�8j���ԜX�h������m�J����5F;e~�Z��c`��#���z�@�p���;��o��������_�سi]a��t�M�3��Hc��>���S��������h��r�������pKJޱ���es�#�\[��M���� .���.�� D���������}�ͭ6�/��������'�կ����������xs��}�;T���xJ:�v*AѲ T�ix���*ӱ&��+~�!
�`1b ����;��'q{s�?s4�T�_��	�Y9.RQp�ߴ��@B� k`��w�'���=�[e�T�+�9�`�rT�J|����*�������q��*�PIYg(.i��y���9���Ɇ���?"�J�+.e�Fv�yԼ X�hE���֣�C�_h�%�*7:�L0�������tk�?�����T~����w� �^#"S��R���׶c�ف��3����'"��|j��٪M����4���!�C^�OQn�O����X�Y��v�:w(��>��z�?��{8dX��&n�d�[��-'鱮����&�;Es���b)
�߹O�+l�?�Q�����wڂ����r����R�����_Ð��YP��_u�Al�w��t�u� ��}��tІNW�5����H[�qٻv�rY1��aT8��yh�2�s|��A��1�W��ŧ��8G��3���uLጊ}?*"�s甍mmn��M!��ʛ��H@R�o�1Fv<"��_%�<�3ެ7�ln?��-�F"�S��F]�H��;�5.��-礒�R�,qڌ�Ŧ�bJ���Z2wn��Z������6�?���?asK�tN�ܑ*�?ax)��9ѓ֢��	9x�/�lucD�7�\֢�O\@l8{�`�i���~����	rh�.j�O�+�~������֛\�G�ڂ&�I[��D�oa?���c~���wS�����[�m��sZ�.�6��)>q��D�Oő9T��"�(n���c��R`<
�0ѱEZv�_�6K��:=}l�.�y�U��	{��?��~}!{�/o��Y�Ý	���E�}ty��^�+I�2����084�FV�P�N%F�=@2wU�"m�i?\�7�	6���%^E���Fkh�	��7� z�?et2Ou�����^զ�5���L��&z:qt"#�����Z�*^���ڐ���}�u���j�"6�s3ouc�on_TH?��6w��?�G��0^��	bg,��շ�O*��,�n׈�Tp|��	iwn5ՙs顉*&��c����<v-���������q�Fڝ��ֻ���V����-Ty+�w~��[,�y�5��<��1�]���gjk/4�|�۬GFrv˺�kJ�z��G!^��P�P�iQ�6����[/s�.�r8!!�|Lj�x���s�>R�%T4��7߈�����'��?����K~����N��*�X�
����J�q�&���Y7z� ���B]�<�7���y�l>-��F�n��O?��ڮ}3d��%&�����	2u�o����T�c�e�'y� k�.��@ξ�����<�'����g�5!���v������GO*�'w>W�{��>9�ӋK1�m]+Uw�m,��F����ߣ�D�z�����G]�s�y��K����f�wH|5���d���V3���߾�m�MbRnofB�X�hYI}�W��;���?[�~��e�I70�b{��9��3>��1-E�~��'/^ڐ����.4��pWE��6[�8�Yw����!��O�X��+ln3g�fk6HLlnkn�,k=~%��U�S�"-������qHL����|��d�ps�D�>8杩Cd�K��~I(����~�7yt�(�a��v�zOdb��b'����Ǵ���Ah��sZ�ױd��]�K>|8*�p��q>��e�4fC�?_ԋ�8���~l��ؙl������y�羮i�����/�捴�C��r��JS�Fqu�>�=ls��:�ʹ}�][黟�߼!��^���H�잴c�T(�q��e=�l������os���?�s��%�X���&8��lŷ�*;���YK]̥!үF��<��ܽ}-?��	�#�X6��s�]*���myF v{������7�}� ��!A��X�>Ops$�+��*ݤ@y&���-�������e�ۋO���\wW� R�v6֘W\��$#������O!�O|le���R��-'�:��W�򨋭!��h9����Ϛw���ղ��fr���'8��BD�K��~��af���T��@�r�=v(���ƅt�f�wH�k?���Ç��V��+{����U���,.��9H�J%�[_ ���3o\A�I�N�������Co>�k<��y���;�g(v��_�y����%�uSsX;Fl伪������oǱb������*o@l��/Z�4e*���	El�h�ZmF�d���Z_��";�BH�l
����7��s�D�7h�ǶU�P�+5OB���[ѪI�s|����5�����{�o�/�y� κ^�A[�t�����/N�v�������N�vg��EZ�Q����6�K��>� hB7�$}ú�nml�F��j�������O��\�~]N�!%��<র��&�kZ����g{��?����w��/�]�#S�Ά ��&p4^��Ñ�Dr��#��l@�	!t��}��\�+~w:��W,��Ed1Y����'<w��p�x���9���j�f�,��%��D˩�����G/X�?=���bd���D��Xk���.�PR�=�pM]|�dMؤ/�����ې�xon�7�\Y��/��J�ف�A�j�g('S�k\\W�ke�jq�\ƶ�y�JTt��F�3��D*_'8�S]�sڱ�@|�?�&�JU�;v}�0�Hq��C���� rl�����5�I�Ig�<X�l;�ܵ��x-�c��኶�V���t;X��:���
�u�}�sh}7wn#�~���%���mb�P�?��+�X��˺X�����OZk-#Z�}q^6��%Rt��kԑ!������!������2|1ߢJ�B����K�1���_M��1>��|�"�z��m�)�s=;���ewp��`U�?���!��Jײ�64���2��5`A��-&�����*��1?98"�9���9'��Z��7�]�P-���q�{�6n��A�ӥ�pl=C�����(f��c���lnݞj; E�kD��{��W�[�5*����'_���\ް��e�f)�p1g�ų(������쓊���B�;����u&J��j_(�ʎ��������@\\�H�N)�X<r�^:���a��W9�[:�<�a>	%�R�Di(~�h/�"ǑM~Q��Kmlǆ�>�(3�mAoTd���i?�,q9����K�c_��E��(9��N�Θ�[Wo�J���W�`�b�]���_��k,,ğG��qA�#�7h���yM����ǚR����}�1��}̗��l��f���o1+$�rɦ���@����Y�σ��
���k<Փ�C����{�nc���t� �R��斲�<&��Z���Y�.Jٞ�?��NE^�BG�K���y�������o!����t\�vֵ̭��h>�ܭ��J;b�O��e3	6����h��ϧHn+l��9���y�K�@֬!h�u�?d�C���uc~ގ%������8��)zmW�������sEv�����~d����޵���Þ��(y�n`�U~E�Q��3��w�w��<�V�C4RWp��׾�@I�aZ�,<Fw�d�/$�Q}?�L-Z7�tkV�g��u�Un�:����uq��=\}~s���7�]z��J<�e�]ƹޛ[nH*��n�5��o+�P�^B���*�F�)�ί�Ԙ	�����?�C5d��$$&�r�ڒ/�y�+�q*���8��n��M��ton���|�F��ogs�����|�������gn���s��'#`A�^-x�͈����έ鏮��Ih���E5y� 0@Ͽx �b�w^����ч&���vQ�k��T�}�F����=��y�c'S�'p���hoxA��xgʦ���f�T�<&f����aQ�ڠ��,<cK^)c�y�x������Ï0x)�;���ɉT�Q���Z6k��bk3w�Fb9�\J�ʤ ;�C�ό邖m�,:́��C SY��|By�����.&=c𕰹�?�������7��n_��d5�!���+mJmk����X�?�ǆc+��<��{
)�̢�r_��r�_6��Mx-�x�97R~�����>�󬟾C�TZb�X��l�.��8�|��dN}�U�%���=�wu��́gBO@Dn;k�M�1ݏn�����ܾ��T��&,�02B�v���l����$=n��~�,9�QO���¦[���i;H~��O�6
����l�u��_8���ga����E��]Ӏq(���w��`�}d��g���'=b<ܹ=��F�oDb���ǐ�+߰Q��W)���x/�|�NY��E��^Mw~��~��w拢�T�����֚���	b1��8�&��/ȓ�k57K���I|�M�aq\���}���H���?e��J_���ֺ���ԝ�_���?���/�����|�L��9ȿ�u��i�i����AzR��'� (u��RgǠ�����*��M4i|�6.o>�ɣrol?�N.����]||�$���u�K�'�l(�]a�C���=�|ǽ�ت�Bb��0���Bon��\h3y����	��D��n�������\X�5�B��"qPp�ݿ��,��J�NO�������w����%�b����M�(D�E�G ���阃S^���!g����3��;㱝�����D�y\�f_��j�M:��] }u����.0罹�A<a�7wF�Ֆ���b��9g�U�y���@G��V٭9;����E��l�zλ=|"ŧk:��w�.��Ƣg�$mT�7�]�������~��ڻnbPl�3�i��oL�G���]~3?��ݍ��1�n\�%�����+{B�V�<�"�}�ɺ���9/8�C��	9��>�b�Q���z��-�aƟ�[�b��_r�Vi~��$HQT,�`���|ų���{U9�g�w�'��A�7'��-v+�U���=͘s%~t�z�W<�O��`�ͳRx�c��p�̏"�OQL�H�|�or���Vg3ʛv�S��w*�O/5/�[�nQ��]M>��?�������m�}�����w������������6�� � �� �[�:�����s}O�*;a�����'��8d}B�p"�X��O�_����9�ou�^��-���Wop�wY�bs2���M��z����+z����7��iXA�{p�@�u0�h�8�w��E�cBZy�����
	��/R�*�'^���6'qTǦ��q�}T%>�ʏ�gbLl�`���u=����o��{�]y�8�<��+RC:v<�L��?���9�����x?Ц|�l���!�h+��z����zm������"�jϳ|�s>?i���s�X[Z.�1fPJA�)=�3�R�HU���8���f�����c��úĦ�6�6!��\�o�~B����]�e7OdO@2[�WP��n�*��o��w F�[r�c�k�y�i%X돲����^��u�<>��~^�F��� ��_��un�Y	`��*�gc�i�fpyu�q�{T��})xg?b!��G�W(��Nn!vj����1��sFl3vS��x^Ϩ�᛿�u$[����:�i�m~�e~2?-��{(�/���c����`��"��ǹ������k>od�u�Z�5G�xф�{�R%����css���;���~ﴹ������C��P�6Nu�y>+0�lf�h���sFe�M>��H�Ջ)>0B,؎��{+Ҧ�;�\���U��M�jb����|�	�#�xC'���Q֗�x������'��c�h_����"Wp�u�;�p�#_��)�v�Q��&(����\�c�jߕ��rד���Qo?�	�)���	J�*�mړĩ��}��G�t{�b"vK��=�����l~ �O���m�����ӊɦ3_�X9��iB�<b�3w�����缿i��7�j�����#�R�tA�0�<��װܹ���^�$�o�����H�uC����ȩ�؊WM��o��7���c^bw�o� ������{G ��z~t�G��ݯŸ��w;�+�:��s�H����CY{���k��?jn�H}���k�p�����P�����\��������%��aqu�P�8�uo�2�N�!��nx�oE��������wP,�f�E�rg<։ù�����`&��)�$��g��'����G�&�����e֠�U��=��/?�'ᮄ�1�����(�ΊOڷ���_���έ'�[�ds.w��ln��������Cfs�P`#p�N&���R�!��1u�B])O�� �N0���Dy����G�f�*.�/^#+�Uc?��O�/:(��sg[>q���<���@�"u�/6����ѓ�w�k�.M�H"��Do�~ԛ�_�y �Fֽ��1jP&9�۟3��R�(.��A�gԢ��WM�}��8����<�8mo���!��g &k�g����c	�/�l�"k�N�]��	���	G7�8��x!����-�W]��Οd�>�l���\S�|��ھ���A��b[�r�2���8�ȳ���6��[Ke��)��Gk��0�5���#�J�i���z������,���ͭ��im�� ��ܳ֩{��3�9�����G&��{�\dn�Ş뻼y���vپ������k< �z;�����;��Jm�죊YR���zr!��豹�;%5ٙ��E�X��h���xA*�t�NB<�q3���V/�1w�GSh�G��I��U�y��!�4��󿜅g�Ę��hC�?/�v���c�R*ɩWy`Ǘsܾk�hN���lVyi�)�ﾹ]K��as���" ��C�����g��mD���,*� ��va�UΨ!5����z�7��ә�[ː.��*���n'J�U旰�=	�-T�Vw�p��� n�O�H,��e��"��q���l1ҭ�t��ǔ�V9�y�Gf���$�Ўkt;Wz�C�Y��m�6�W����`�l�a|��\�ob�����!�\T>�X�jK�ϥyN��xw/��1�ZL�㰅�Ƣ���} w_tw��Q�6H��X��lN[�uȯQ��-��ƶ(��g����$�����q�W��<#Y �%� 7�X�S������y:�NrB;����2��zG\�J��W��QVɩN!�|��H;־Y�]\�b3o��O��P�aEöJ��Å7���҄z'Z^�����.T���<�M��+�P����&���I�	Rfί�0m	;���"?ֻ����-I}��K�����R>�C�_�`o*��Y��|Y�9��]kL��m�{������~S�1@.f��G}eOȾ�zE`��ox6S��V<�O�ݡ�W��<��|��ѯ���gVq�pF�����lͥ�]��[𦦘�p�Ж_��ql��R�������b%uś���\U2Xj�F�z�~�C,�ERZ��Iʴ��/*�#6^�>q�z����s�!�7�.L�=�[mqr>e��g����Ɍ���'[e��z䋬5�����f�'�B�On��Aż�-��(��8ʠmf�E���#��v�^���$c�B��E���ȱ��M,����֜�i1kQJ[G7����ʂT�,�C]r�����̟6��[.:|<���n�����ؾ�:�Υc|f8�8�����S}�Z�הv�t������=�x�&��E��yf�,R>�o[���Y�跈�@=�)Z���sg�Wc����n�$+�$����Oż�>7��FN�vb�K�ix��M���:V����*-}[�g�7ɬ��9����H0�Z�+����͹�A��n����v>�3YY�\�*�����^�\��!��Y��Qm��;�����g�[*#\^�Ѿ��6:?�B�O������>r���d����P�<�̫~�S�c��vPf,�{�z|�_y����{|�;�z|�_{���6���4bŃL<Q�B{8qpP3��Ԉ�fh�<I�+�w�v�pZ��2�~�u8i�Y��杯	PUS��2�(p�1Y�2���������M���
�/��%��'="Nw�ќ)g���s�β��1uޯ]}0��8�_~��^	9Yx�سN����G�Ba<��l_^XIJ.%��Nko@�Y祪�<'��?Ν�p_$Z7dN���:~0��0l��yE�X�ZD'�U����;,��J:��;�IMHJ���\k	�uj[$�+��9I�<G�R%����;��/�ð���j�r��Z�p�ǩT�~�,T�_j�E��]`X��ט���8g�u٩��:h��vb5VXUg�� ��cCux7H/���羹���>�}���u�n�t�]����tJ�#.�'��)l�~(*��ԙ-�K��Cs�q��[�H]n��m��>������ޢ����U�ɼ 
�4�+��|��X?V�Wڠ[�s��d�w.��������4�[��5|B仨u�[Ⱥ�����wkY�2.�횚�z�d�1�.��Ɔ�����o��.��G�S���@<֩> k�ĉ�x^Hi�]ds�����~ۛ�����k?s˃�.lN�"�5������p%7����a��ϔ��<�@����¼4+��)}*�GR���B͔p�E� ���Y~�םD�OJ��~i˗��'u�'����q�d�����wRp�� ��Q�����K�
[*{�b�V�v��A�\L+5�`�.L8�6�T�25�sƐ	��)��MH�/+�@V��#?c��s��ñ��*+	2�����cE��(�1�!m�ukި���{�^�?Ŀ�~�����d��NX�<ӧ�ПX��-�voN��Ӈ��%<-�,��3H-���]��O�e����tP��������~,�?"d����ȫ�^��s�H8��n�K����:F�~����h*N�}��/8O�������C�r�ē�Ǚ���W����3k��qtuN��<���=�m��tB��m�x,9aV;l���D�?���3�-�-��x��#ـ*~W��Կ�����P9�x���ҟe�}�νq�=@�U���cr�����'�A��pc^���u{�H�'�q�r����]&)�=G��hD:�n���d�ɂ�^W���-��/_���%_�;�1>�We_��F�E��flq�"8�6����Zx���:�=G�!d��Z)�]����g��P�W�g~�����?��m��'��C���5���w�m�X�/���i�8�A����3����S��QŁ���d���<�P���ٓ��?��l�H����Ƙ\���	�.�6�]�I񑖬S�Q7�ye�^yl٦�b�tB�;ԫ?E���4u�Q�פq��G�n���~tR�;*R��K�(�kU��A*&O(W��O�Nmm��*�4�P��!���`��B%S�G���'���u����T�Xr�=�i�ůl�;뻗e���g������{����+Q��Qb^�b�y1}�8cD�״�e�6��A���~-ZV���|�Z�#	؎�U�=�`�{.0�����%rׇc8n�!�E*�\6�)��O�*e8�Qv�'�RKZ�Ѿ������hB��А
ȏ����:1:]��62m�X��]�7�g�G��fx\a��
؉8s`���+���K6Cؽ!���ᚶ��@���D�O��~C��1�yze}J�PW�G	7��3�+O&����}�+�n֩s�6$g'U�cw��I�lb��3�%����D~{��g��#�X~]k�7�Pl⧩=��}"�-�Nښ�Wl���f����-e�L?�Io|Q�'k�ڦ�:k7��x����׿�[�������ۏo|�s�F�	;emn�Y���A���0Ly� QS�+�-��|�W�鉼�` �Pw)��v� �m����B"�~��A�w,֥±JA�>���ڒ�E�쑐�/D���U~��/)�`��\\��vI�?�fy�c�vُ����̢��A;��Qb/���Ł���-,��h���(��B�	�TF/}�,<T6v q*�k�bTPe�-���b�� v8a�D��j�>3N���"���>j����"Ty���ǟ��3Z�-j�h��}�������s���1��tJL���OV{�p�V�Y����-+��:@�&iK�k�/6��<LUf3#�-"ʜӬ�� �)lt�]�W���0U�p����TΠ��χ$P1M��WlSNrō>���wO��w[}����h�k�A���q����^p���>s�&�x�eH+���
��2~U8���&⌳�Ɔ��˨ˏ_�F!�o���=Y����M5�Ϲ��wF�k�p�ݺ���<�����g}?�w��0�6f]p,���c�O>���)��)��dc�}�7�e����4]�*H,����Y��K���f�=��6�;�x�/���U��uS|��u��h���ZU|9�7�W��O�}�ۏ�������������|,���B��2�M(7�%�؂.�Q�8	��Ot+s���_�b��E>1<�l4_��o�'-)r��.�M��i��
@o7����.�	P�ԗ� &.�J����EN­{�D���Wn���$��2s���*��9C
t�[Pq��:�3�䜴<�Ņvt?��v��]oj�-��"�y�c�ln3ߒ70dR��[(�`��U:$���na��[����!��,���]�6�s~=|Z����x�O�ڿgM�����D����>���v�a�����p�O}�Q�I`=�?j}������k��h�M٩d�������X|�V�\�H�~���w��dq�S�~�[ؤX���۰�~�α��
f��@-���o,���k�dUe��;�ω�mdO�Rl�?�^s�>7o�=�<7g��Y^eK��b2�G��Q^�b7s�d� �π��c��uS�{�q}n�T��O{����t#Umߵ�v)q�@"[E���d#�y�{k�dgTXW��y��/���b���o��ьF]�Yo��	)>�l��b�pƙUe��ͭt}GZu�6�~,A���7�����wn�m`�Z��b>����iE�xrG���N�ƖŸxw8�\:�X,��:��73I�n��ǀ���Y�m�)��"qt,�ޗc���(%�!���Xx��?��n��c��QV|�AO�H�H�	�8ڹ�P���E)ٻ�g���h��N�1����0�fƴ���EJ2`�b�eQYC�c8�U�<��S�4�U'�$���p�I��.>p���8e�Fx�U��ew��$�MϔS�1�?*���T��9AV���u`'�n�⌜�?��;�1���j���d�U�������%4�c��y�vu�C�A�vd��L��ǯ���Ni�t�fR��(O(/I�Omn��^縰����E��l9�U��K� ���C���4�æ���*P�s���r��lv<cx'�$6��T��2��6<�J������*Lꕞ�6~ Ƽ1]ᰟĎ۬?U�=�t��g|J�Ǚ���U��V���߹��b��Xw���� ��G�,�ۙU8�󷮇Wd��cBA��T�/�Xc���/Sy���1����!�#��#��cc�:fҦ�וK�C��U�%�<�m=���Ue��G���7
ِ[�����Eon���_��fs;6ت��_�0+�B����l���sĠsb���^��&.��#�B���.�"�X:_�Qi,\H�O(ex�M/o~(�8�H�w :��D����L�n���D�#$��{R����Yb��M~(*N��&�2���n>�!�ll��463&ԇ�.v$>i|�U�ؾ�J��Z���P�H8-y۰i�엞��s��ذG5|�>Cœ��W�T׽/�ճz�\��~�ͧ~�u�5�Z�Z���}���@���9�y�������o�ί`�N��g���}�sv�.�E������!�^c|#��[�~���87ͬ$%&=�}qפ~Vl�;���M�S%1��_|QH2@���Ia5"�G��Rڏ������C���Xf�2�{d�W�����ހt������C�m�T�&dk�I��v��0�����X
W�g�.olX�C駯�H���k��?z�ͭ��;�_���o��ه���'�n��΁����.�~"�hH�^�s?��������<��[�roh����k�è�t�H�t��T��c�K�:�s>$�۲����jT�6�6������s[��?���%��6'z4���Ug١X�&gE�e(Ζ�z�;�B� [���0c�m�7���	ۮ4�Ⱥ���.^8ՙ�:
jCΒ�7�¶i&�-���:�H�O��F���)�>����6�r8�I��b&�m��9զ�F�k{�������~U����S��]���1n���lTH���y��/��۲�p��z� ��wY�,18��@��q����\�;l�NU>݆-�O����@AcG����A}e/��%sЯꏌO7�ր�.�^ņ̦O8��;a�f#!�m���5n��ll�����;˹��Q���I��Ab�\��N{-�;8�u��wZ_�B�3���vYÇ�	���U@\w���}������b�n�x|<7���g,����f�W�n1���_���i��VB!10Y/{��ظ����Y�K�X��mm����Dp�m��������S�m���ߢ����(84���x�O�� ;����g�Jq�U����G���O��c�O���vܩe��R���-��͸]���+��K���V4&��5�dG~���mn����_�c��L�G�'�����������h	��c��b� 9߭�Ά	� 䂠��7l-&f1�M�����j�+凼�v�n�����U�I�)H{��D�g~��~�.��5$�6l���EL~]�C��TR�vy�[�]��[���ND_@*��P��ױ������q���IH`3�����uچX���]�oD�EGV�91��DǊ�m������ x�&�y�1ί�8�	7���O�n�x�v�y|�������"�J��}_�%x�JǺ}|�,��֙���iQ70ou. M��s�)�[Q���������
qGE���26�}a��Jon_]7��nڟp��-g[�\�q��U�(���!�_�[���p�*����k�-�)O}�3�"�('�C;N#��ָs�0�}� �h��.�O(M0���g����>i���6�z���R�5��\���/w��i����~ڒ�-�������v@|2r�v��� z�����O�+�H�H�s�uG��ld�e�	ao1XYm���V��7��|u��N(A��{ �`t��:�|��̭���G�����2?s�W�)���@�ۿ��ݗ�K�m��@1F&Q�/��-|�s������˃a����Q�%���+�X��K��1�B/�-XTc�(��JK��B��N�G����������|d�B*I/p���
-���I���8nl�es�����*'Ag%�_8C��?'{~�{(QF�F������#M��DUp�8/��TJ,�A�;A��s���0���y�w������g���>��=o!�림 �o����n�p���{�n/q��s����c�(�:�V���\b�*����l���
qU�切���pa��Cplˋ���+��c�����a�5c�;�a�8e~�o�sL����6�!���~�T��m2^}�u5�:��0w��\���9���?Rk����Qa�[3���`\�6����G�A�ޡ�wf�5�)R9ם�w���c����x�2�4_?>(g�t�����)n�s`�� j^_Q���n`UѰ�yR֖�����Zc�E@uT[���������E֙\;B�M�V�Bgϩ�q��	��{� �W��x�46�����<s��o=�ʛ۟>~���<^���������E }X	ia^�X��:)\h�Aŉ����T����0d��/uQ�;����uDV+j8�C���x����{���AtY����@'�oR��
���!G��9˹d��� /1��d �ܣ�&� ݒ32��y;;�䓁����$�"��K�������B��A)���n��<U�ce�Պ�" ��^J�V�@��N��E��O��]�z�Y����S��~0;;`�m�O�Wd�	�'0R����"W���X,��M���?�s�io��Ts��_����[�[ǔ],��+ ?��\�����t�/�"`�d�X5>8�t^��j6�o^�����܊j�y"H}�Jg�p�*�|�W����u�]d����apK���g���ҽ�oO�:/7b�}nn񃫴�/�j�3��#oc�>վ;uU��;������>�g����ܐ�,���+��L߇�����"�:#��}x�F$C��8��1�VCD��$M��K��[�&�V�����<�^�jt�>���kgh>���1?HW���V4��/�ɍMon�|���8}ݬ;��on�|�x������ۿ�S߹�c	��-���Q�c��=�iU��^����<6�I�t8� �ؼ�^$=v�|k���]�4|�5�M�g-�o��c�ud���n 1�B#�#�ÃY����5Nw~��;�k;w ��:�1�t�c>��	|AG�n&����;��"�)���b�5W��yө�Ŏ�Mğ�9W5Я�T��mT���2��? ���4��v��T_������~�KA���@��խ���]#{�]L�(}�%ɝ� )�W!��&��@:eת�pyA�i�m�]֐ϘaǩЩ��C��eI�z��Ouo�/��?Y/fl���r���7�dZ�I���ao .r�_�Wt�ҳ�w���v��q<;/:~�1v�~�7@7���>!��V���c��[8��gA<�쎍��}q�t�)���m�9=���ʍvm�	�ו�/��8n���K�]j���m���Y|�o�l���r+Y��Ӹ~X��]-9�Q-��úG;���e���V�hk<�;��f���.w5�@��6��?VҼ#�[����J����mI&��[�-�]��8ʠ;=�* �Q�Xi�0�-`^��w��1�ͭ?Z/�h0O��P�N�2'�����l�x�����hƥ�X�����L��k��Y�'�n�O�6_>*^�9�r2�*�	U?��$��x���؅�z����E����~N�'��@{􅡔��e�)�>�{8d�q��[|&���� ����9�8_D=�KA�+�ad��ﱟ'Ҏ�k��?<������$�R�Y�g���B�)^ 1���KI�9���υ�9QuRp�<��Re�'<�b*�q��؈.,�2UK���[�s�7�;�l��O��wFl[H׮}��w��^�������Yx?_����]�vH]� ȸ'���.@�H�}�*��1s����6�A��\��Q�}��>��X^6cp~i��t�;ǾܐUǉ	������o��y��r�[�����<�!�3?�,��n��q}�*�*e��j�%��?+i�̮&Ձ�����w6�ئ���]K���?{��~z���;RN����+�D<d��[�O���i+rS[ĝS�"�t��]c'�]'��	�f�ZP~��#dnM��Uٓ9|C��Y1�hy�+{L�[�j_��7��4O���;Ԋ�U��P���M�W��:FOP�$��gF����������_��HcC�Q��;�ESPiD����_��'=���m����C�����|x�ǻ�X��>@Zݠ1.G�z�kX\<j.�O⿏���|*i��7l�^���*��gh�V�.�8qn��U	C��7�i�k�Ȩ�)|�(�D�u�؛/�H�	Q@�hN�d����݈�G��Uo�g�����$Vq�_�:;����+�mж��+��/n��^6�C�sLW?XH�a �� ߕ=��D���N�y���ڌ�6	Cw�M��nm1w��/l�'D�q��-�'��U�<������c������t҂���ٿ��t݋��c}���㔗Sr.�&lf�%Y�S{>���^����w�߹=ln�s������
�+��Դ4�h�4^&F�S�����A�zwV�����ӡ�S卭E.���n+��M�K���7��y��Pyl.��q��	�0��NHTȘ�@Tzc�jB��8b�� ??���/2�N��Wf�L�.V&x���!��&-[���P}0.�mR���}��|�TDJb�����!|���?d��FN�{xG��9���w��N���gu=.w-D7�ug#:O#b���^o�vH��<�F�p����6t$��R��66!e�h�f�M/r�p�������䏋�	*��伃Ĕ>v-�M
��F�C:��h�>ud-�t����K�;Ӣn����n@�}?Ѿ���~e]����ei��b���j�/��^����e�/�qyv�.h�O���&���܂E�����wjNb�ɭ]1e�>���������1�_���Uq��Tz�le:�,�!
��lEާ��!�7֗�Rd���~�k��ORl��'�7�dʵ��7���i��N�I��8��u�:K�������esKL�,�t���ln���ȝ�esKc�ݤ���i�8J�)u#�)��s��!�C��'�v#�3t*wo�Y#,�:��S[��$�-��dn;���t�ɘw�ys~}U�m�h��Ɩ6��e�����~Zڴ���i|�U���ձ��q����m���[fcI��qGn���W�WWZ��{���$ʦ`�`�S*�|�c���L��n+���	:$6���޳��_��<�����T-�t76���ڶ�����HM�K|��mgMyYȪ�u��;;4u�;��ls؜Z&�{ӛU�L����������/?�7����Ŀ�-^��܎yHQ;��C�+'�޼V*9Ho�B{6�����ʍ*[�~�k�߅P�c��Ǥ(��7�̩'B��v\L4��vj������:t�{��Nx�Ŝ�[�bbGt�C���O��I}�OtuN��6:�-�TY�hŝ"��Ȣ�7����%��ͭR�~?�7����P]{�~h�llGW*�y^�k���<6��� ��5���v���H9�r��:L|�k	�����s���g��ۏ��VT|��J��X�0ސqc�� ��E�.�#b��c厯E��z@R&������� �G�#wЭvd�-�E��֭��Ug=|QM�wh�FxRV�Y�k�^I@nUӡ�;(9a�Of�O\�^�鰸ϫ9_mJ[�n}�����%��M��gdFeQ��͎�"��q��3�܆��V�W��ڞ�TIj�;��M���6jx|חlN����� P���z�U1��yn��TJ��@tt���::��*{��k�'`\t�W�?�]��"fRA|2֖��j�i6kϚ��m0dV!�X�0	ΤԳ�յ��cޤ����3��[�X��h�,/���L`�_��#�
Z��?:�3�F�Πq�z[���t�X�[�{��wC��H�+�\vYB[,1��j2�'����{O���M�������jC}�LR��W�}-���x�/y���I��hW�8����Z�1�|n;�b��6��@mƱ=vBp��J�$i��J�B΋7��K麮O�����|�F鋿��VG�oK�I�ve�A�l:�c`t0�I+T�	A�P�;q��:������պlt��Sˠ��H>�չ-纐��ߐ����Ыd�����{���n�Tj[A�3XAɫ8���AV�ق���%���'F��K�l�\J}O��p��4�rj{=>��N
d�vH�!Wˀ�Lz�i�W䝔l�M,��M�R��J���w�o�/�+��9�M��5ƆX6����.���Cߜ�ӟUX�����}�}BD�
�}��k��ia�ٯ��IQ�*Jij�x����q�f��!�:���2�*	*����_@xp��g�4�|�F�����g��1]���/�����5Y������%�P)�ˢe����q����m�mm�� ���gۭc�θx�Y��OPr{�RUӅW����+q)�n��-�x��Xi��$mƙis�b[����/ܠmp�mu*8�
�����ھ#2y��X���g�M�U����ݝ��V*�c�~��9��	�=��gΟ�@�G�k�^�k��bw4�Y�*h֍���cc]�iln����p\�e��T~d���y�<�i�׫*�Q����|���/>{���׏���7�՟����?������{���_��v*|�O��������ds������L�u����4?8B�,�AgH��O\�6ؠ�C��A�\�*>a��-�g�s�p�l�rL烽ƊE����U���f�\1������^�~�c.�����CD���|�Y��30����Â�m�b��v[?i�`�g�O�w�#��p铲9!�'�;pn�?��:?.v������n���`7�w8�^�,]�>��]��&�q�����Yݵf"��۠��	��t�08�9���P^x��OZt��`[�v:�����栊{������c��l]��c	�_��1хK<R�s��Xëp\NA2�����K���8���Oݽ�[Pj��ž��a��nT��Ψ��>�A�|Qg����z3�����7�wYz�"n�g9o ͱ��f���G�~�P��s��b%��?�};ޅs}�+0_�3��J3��\��7��G)BDK��TI��(,�D�]8U���b���D\y�-H���X��w�>���
�����X�;��>Y��%hc���k?��	����O���?���{��G?x��������j�'����P���P6��&����M��F�ą����������|Ý[���r'ckKni�5��FG�24���@g:mݓ������E�ڕ)ocTK�jQ��>2��q�����1�m!�z����8�Q�d������s�+��%�CZ1-����=�+$1ad��BZ�g�x��'�c�|�}���������±�����b��K�~�2������+��T4D�m^�-dC�_�T��Z�ڏ�W��
������!��-e�qq�������V˲��Oߩ�M����[]�d����>�,?�X.\_�@~?�~sA�_�#ϔ'�a�e�	��It�w����!��>�y�oտ郕�����|�Y7�u}}�]�r^���Sd��,m�l��s�C�1e��N�?�^����(+u��Q$��]��b=6�J������j��%�ю$g��6��=>�"��wv5q �Wv̶�5_�Z"�ɛZ6۬���.���ɀ0��py��'����<^.�Ur��v�3��긁�]��S`|�Lo��|�;��ln�����w�͗/>��	��X6��㪀d޾�?�ܞ<;N�n�
C5� �l�Op�b�p7P�eg�tg?�z���k?����oЭ���Ҹi����1�"�c$�v��͙^�c��>�XC���>�����]sf ��!$�cJ�A�k���]K�Ԓ�5��������Fb[� @&���ŏ6�"�C�{s����_�\>6[�/�fFU�*]�G7�����E��s��քx���]sTg�WN��2���PR*�U�3��B�����y� k�|��/5�lH�ɒ��?����c�����K!�v�$�q�ܶ��7_@l]����(C�Vqϐ�z�E5���������9��u���=i[Ò>v|1nb�tު:�����z#����3�_���6bנ�>#8�mX�F�2��o]��y0�b�y��K1V/*gc�]����3��IP&� �i'���)ig6�lz���s��Ȱ��܄\������/��ˇ�y�R�[�`����_o6�N�⍺!��Xd:X��#]�4瑤^��e}������ϵ���6���ß�������~��p�6�`T'vcx��C"�a���x\(�f�+���\UU	�������./8L�a�-P��R�;�#�gO��Ļ��}dy;Zs�Aw�b�X��k|Io���+c<7��W:l_�v�As�ڮs�&���H#DU<�&�YLu6�Z�=Hn�����H�bg7����I��^��_1u��+v�}���.8��B7��K�]*�樞�l��q�*o�%?tV�ʻX<t��>�֢o��5�Jc�-��Q�\L;%����z��=R�_�*�<㮭��*��ͳ��)>�9"��w�܉Ʌj>s+��<�M��6W�#0�8�|���c�S�|+�v�c�c���v��� >�.����(�����'��I�~��7��h�$+l��*���*��{�ܮ�/��`�8��o����q��\�;��Y'G��.���94��%���NI61{i�Թmw���2g��g�:3g���n�A���yPk�IBg�gA��(��Z�y��]6�0�N]*��y�|�e��C6����Ror_)����������������Ǐ�cs+9����T�yeFj�E�Kr]�9Ƀ�pl�N�e��>��c��ŷ�j#��h�XT�� ��&
��/�:tL�Ar� �����Z��e{"���jjt�K�誮�83K��P�X,���H�E���dH{�FXѡd$���T�a@m��q������汄�q��F�Illnw��g(;���N-��PY��{��Q1`\C�"du�w���bX\�DW�L۞�+=��
�������p��0�S��4Ť%ռT���|mv�9���ǒ1�����D��G����67'�hEe����nN�[P��v�0�J�Rb�m�FVv�n Z}1�8��'�6H������_��Y�A���-����ʳ�-�F�b��Wpe)�ܬ�@���o�vv U�]�pB��M�˰=C�sr�;��{�_ۈ�s�U��s��F���?��w?����6���W��^�ݰ��9�ˎk�0�}���xө?�s��k��{/�|=�s���\�c?�?���e���+����w�����~mn�����~�ߑ��S)Jۋ���tL/��k:5���\�9v��Y�ٌ��ѵ�Ν�f�&΢=�s"<�%J��T�.�H�:�V8��ZTg�wZm<.Ю�x����9�k���;�b}S�0;u>n�⋹;9������֓�"�c�i�=�=ح9���!G}e�d��mZ�0��$$�sD�g���I�v�9W���X�t���>sў*綄?jIm��W��.Rh2�����q��{�m��)����l�i�;�7���+=SoBu>dS�_4�9�M-o$��ز,wv���ˋ��6��\���G؊��v��d���`�x��uS�$���������5�S�3Xu��-J�p72��B���S��tL�0�O?�bʸ����VVw��Z:��y�`)^�_�9e4�V<ۣ^��a��M�6����,�N(o>޹}����)��p��}bʎ~8�4J����Ua����Ț���XD����8K�����tt����!�-�>H��!�[��s��	�7�����B��?��O?��/�����%�����&������'h�Qj��Ȣ�CfN�Z,K}=y�_��y�?N���RUq�P:Ga��T.�T8-���� X�Z�XĻ������_^(; ]��{�M>~*�����X?�(�Ő?�)�܎n�:zĝ��e�.bS�]Ṋ<�v����u%��!]|���E4�q*�a��d���s�q��c��eS�BG��,ot�W�+gJ'�7�]�N��k�@\�Pe�ڃ�T̘�`E
'w*d[�������v#6P�A�+_�f�M+2�c
�)��2������.>�n���ڶ���zl�sSe���	�[
��!uo��x⫬�X�X�u�PO1�Cl��:Ӕ���� �n����C����k�(�aS�b2�=��k�^�d��?�ۼ�T�ؾ	�H��zc��Y�kMc�N�����,��j�X����t���b�տ�K�E���aڭ�Q>���|���߆��q�.���u�����Q��a��xQ 6�r`���}~TAɕ��(���
Y�2�/D/���ś�w����������ޏ?��/��_����a�b�M��G+��gd�P����Y#_R��/-Ҿ	�lμ���z��폍�o�,�0Ά̹#R�(��f:O����7���Yv$f�׺#ʏ���Bg]�CL�`V|��E���o�cc��ή�ߠ�>���}��@j��ͫ�z�l���1�F�����o^�P(�M��^^�X�D�Rx�Tڄ���C�R� ���b�N~(��ӎ�'�:N��/�m��1�����菝=��4��l��ƔWn��Zp(�<�t�;ul�}
c�B_������P��N��:.2�J����(�i#v�_�#��t�b^�|�Q9�A�OT0�pc�����St���D#���b ���Ҡm��2+lm�'��Ҟ38��œ���2�ŗ���Y���H��
S�3�In}w��{^c����?��Ty��,U�V�����G�iE��X�>���F���4�?}"�b��Nds	[�s�����ũt��W{��7���O�x�b�qs2�opn7]>�ٶT�N�o�C���npK��S��\0i��s����a�.�Q��n{�B�#���Z�j�i�B��y2���k����A��8���c2��k�������|���;����'?|���������������eBfQ�sjOͲc��W�^|e9��W�-�ŗ r�aru�7�(�ͭM�9�:��a;��ˆ�}��Qt�R�����v�� ,W��d*=����6�J=��&@�<���>���[qR����/��?:��������K��/~����"��\8����F��c��_���d�9��i��ߙyt���g�/�e3�����; �N�;�斶���ܙ�[b�Z�IWؤY��̂�5@��=��/��o2V6����
ҁW���G�/�ᡟ�?�r��X��ల����M�+�ϛ��[7c^�Ure� �~)��]69k̎�\.H<7
��E��26wm��ըx|N��;X��+�ue���;�����E�C��,�˿�c���U'�����=ԓI=�Жd|4J|�C�xݦnK�-��?��-�>6Rl��;]�`W����A\}C������|d#����ϱ���ʐ��Ҡ���X!�Qf˲px�����;;��8�$X�1�X�6<s��r6�6���\�c���|��WU�쯕��������> ���D�봹T���x��}�~���ס6p��v�kJV!������m��_�#���۷�?bs�M��ͻ�oOo���x��~����7����v��_?�[���M�_ha������H�S����s��ps������Ӎ-@׋��/^G�WJ�=��,Ǧ�jR6�E������6�,�t���ܷ�"X��Tar��g����C}��'?���o�{�79Ǝ���G�aeMR^�76��9�� *�������xm\���ױ�m�DhR�4/U�u�v�qŮ�$dN1V��H�>���g�-���ڃ8ӓ��u�g�%��!P��WL��,�yR��׵�կ��c�s�y����� Nl\�aλA�6���(
W:����'7�����v������0�����'��G6���k�u ,���ܢ�����h�PO(������ˑ���hZ��S���{�3����Y�yq��> c3�c\pmʵ(1�Qm�e'8V)����/�_�'�T�GEW��8t��e8�GR�� �&�p(�X�'Y'$s�A>u����q�A<����$L��C#u5^#��������O�6(9��@�*�P�s��x���V�On�'SA�X�k;�O�}�ܶT`�S�]��-�M�˻��%�6�w_|���/��y�����{q���ٛ	mU����:��ż�z:f���(.Я��q�l������Qeg��������n*��8D�HI���՘�5���:��f[t�M���^�c���m���_�eRcٞ���_����Ws�����4T���ķz� M±�S��E߂s��4t����_�0���3n�/�Z�L�����p{���5Az_�>��Ƴ>Tk��$�a~�*.C�s����H�8p59��@���Z��Eu����lu�,uF��r�uz��1��76���j]��(/�7�����.�����bꅼmn�]����Q?~�WG�c�������9�Kr�;��qk�� c� '�柤:�Ox�{�g���~H6xj�Rd[YO��e�L����������S�� ����Ж������Jv(�b�k��,q ��5�������b���a�֌���B���k�s}�U�Z�f���X��p���9(v�9'&���u)u��ĪՃTE(�<��6J�/zs�׫���qs���.��l�gO?������n��6�o�����������UZ��W�;h�"��4��[7YymQ�e������g:�D���3�Z����v\-�@�����������B��|#`3�2t��#P�mV�ܙĹ_߼r<mER�g�����ч������X�'��p���O�U��ε��
�R���|�ӥ��Κ�}���\�����6�_R�a�'���׊�yl�!g|un�g�'��Ї2v3�g�������1�uي��g}�ϰy4JI�v��1~j�?~�pT��	�1�o�XU,we�6��W�m"m�*5���"�qF�W��,�����ڈ�g���w������}�u�3�R����:P��"�����0���G�·-��I�̐n�׌�r*^�'�t}�YQ��K<�N?)4�v��[��>���k���ߡb�.v�U�56M��,�)!\��Uc}�2������Su��� �u ��A�������(�~ppX�1tm�p��)J'�;`�ه���{C!�sd(�🥓D����YcĹd�p7��ux���v���u�ڎ��Nh`1\?�ϧ6�o����<blp�~��
/�1
|�<��fs�>�O��7�/�������>�^<���{��~��6�o��~�������FWͻ����#b����&�7cܐ����2�l��哎�gs[�C�x)�]�����&��yT��/:M�c��"�SD.���l;.y CA���?Ci�L��`��4v�oܼ�ɍ,���R���Q����ڿo��ȋQ�����\"��{�L2��V���LM���.쒋��<.�3�9&��o��퀹5]��/17����a��F���d-7�c<� ��u��-bW+e�����uɺ�5w:�Ƒ�@zV�V&�O����$��}���m�;M`��m�):�H���b'k}M���U �\�25��:l�=75�"Q/ـ�kQ��/Q����E=�O��Z[c�7�����%�m��}��vȇ��y8.'j��m�5�����o})�nMO�%�O�c�'#�@嘎�p�<�u��iK��5Ya��c����G�f}�r�е��l��W�H��Ӽ���>��6O�n�h4��1h��������%��j���/��z�fkrEq��Qu��������������ux��)�b��8�r��hp�9�^��'t�b;$�I�#�cPCk6�c?{BotU���vĀ�CLQ�*!�c���[�=_ȃT�b=6��R�H�v��'��>��x�}���޼����'�"��M    IEND�B`�PK   x#Xb�qۗ  �     jsons/user_defined.json��QO�0ǿ���A�Ph�fF4�lSP_�b:m�Zl�eY��E$n�������n�mE�4�ʗ����O*\۱]���W����yw|̳��M���J�B��g5}r����Eߢ�1`����H��C���X��������1����Z6��BDU.YU�u��X~��]�7]W1� ���:b�*��T��G�^��.����Ab���A�0����F[�q�֒i}m�$Ō�+�*$�&n���ٮ3\��x�.��?6[f�Ԕ��[Ў��}����Xe�:%DW��'�Z��~f�4Dx}��4����� ��!t:�!N��	� �,��<=@�Kg�����@^x)����h���x8��z�[�%EEe��'��\�W�]�_PK
   x#X�i%X,  X�                  cirkitFile.jsonPK
   0�"X�l��z� S� /             �,  images/02fd9929-a358-4090-8e7d-8cad28564328.pngPK
   x#Xb�qۗ  �               L� jsons/user_defined.jsonPK      �   �   